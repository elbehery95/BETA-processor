`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Abdelrahman Elbehery
//
// Create Date:   00:31:14 02/11/2017
// Design Name:   BETA_TOP
// Module Name:   F:/Self learning/FPGA/Projects/BETA_ISE/TB_BETA.v
// Project Name:  BETA_ISE
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: BETA_TOP
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module TB_BETA;

  reg CLK=0;
  integer weAreOk=1;

  task PRINT;
    input integer CN;
    input [31:0] IA;
    input [31:0] ExIA;
    input [31:0] ID;
    input [31:0] ExID;
    input [31:0] MA;
    input [31:0] ExMA;
  input MOE;
  input ExMOE;
  input MWR;
  input ExMWR;
    input [31:0] MRD;
    input [31:0] ExMRD;
    input [31:0] MWD;
    input [31:0] ExMWD;
    if( IA!=ExIA | ID!=ExID | MA!=ExMA | MOE!=ExMOE | MWR!=ExMWR | MRD!=ExMRD | MWD!=ExMWD ) begin
    $display("Error in case: %d\nIA: %b\nExpected: %b\nID: %b\nExpected: %b\nMA: %b\nExpected: %b\nMOE: %b\nExpected: %b\nMWR: %b\nExpected: %b\nMRD: %b\nExpected: %b\nMWD: %b\nExpected: %b\n",CN,IA,ExIA,ID,ExID,MA,ExMA,MOE,ExMOE,MWR,ExMWR,MRD,ExMRD,MWD,ExMWD);
    weAreOk=0;
    end
  endtask

  reg  RESET = 0;
  reg  IRQ;
  wire [31:0] IA;
  wire [31:0] ID;
  wire [31:0] MA;
  wire  MOE;
  wire  MWR;
  wire [31:0] MRD;
  wire [31:0] MWD;

  BETA_TOP uut(.CLK(CLK),.RESET(RESET),.IRQ(IRQ),.IA(IA),.ID(ID),.MA(MA),.MOE(MOE),.MWR(MWR),.MRD(MRD),.MWD(MWD));


//always #5 CLK=~CLK;
//always #1 if($time==10000) $finish();

initial begin
  //CASE: 1
  RESET=1'b1;
  IRQ=1'b0;
  #1;PRINT(1,IA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,ID,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 2
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(2,IA,32'b10000000000000000000000000000000,ID,32'b01110011110111110000000000001010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 3
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(3,IA,32'b10000000000000000000000000101100,ID,32'b01110011111111110000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 4
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(4,IA,32'b10000000000000000000000000111000,ID,32'b11010000000111110000000000000000,MA,32'b00000000000000000000000000000001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 5
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(5,IA,32'b10000000000000000000000000111100,ID,32'b01110111111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 6
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(6,IA,32'b10000000000000000000000001001000,ID,32'b11011000000111110000000000000000,MA,32'b00000000000000000000000000000001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 7
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(7,IA,32'b10000000000000000000000001001100,ID,32'b01110111111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 8
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(8,IA,32'b10000000000000000000000001011000,ID,32'b11010100000111110000000000000001,MA,32'b00000000000000000000000000000001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 9
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(9,IA,32'b10000000000000000000000001011100,ID,32'b01110111111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 10
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(10,IA,32'b10000000000000000000000001101000,ID,32'b11010000000111111111111111111111,MA,32'b00000000000000000000000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 11
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(11,IA,32'b10000000000000000000000001101100,ID,32'b01110011111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 12
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(12,IA,32'b10000000000000000000000001111000,ID,32'b11011000000111111111111111111111,MA,32'b00000000000000000000000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 13
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(13,IA,32'b10000000000000000000000001111100,ID,32'b01110011111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 14
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(14,IA,32'b10000000000000000000000010001000,ID,32'b11010100000111111111111111111111,MA,32'b00000000000000000000000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 15
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(15,IA,32'b10000000000000000000000010001100,ID,32'b01110011111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 16
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(16,IA,32'b10000000000000000000000010011000,ID,32'b11000000001111110000000000000001,MA,32'b00000000000000000000000000000001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 17
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(17,IA,32'b10000000000000000000000010011100,ID,32'b11110000001000010000000000011111,MA,32'b10000000000000000000000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 18
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(18,IA,32'b10000000000000000000000010100000,ID,32'b11000100010000010000000000000001,MA,32'b01111111111111111111111111111111,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 19
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(19,IA,32'b10000000000000000000000010100100,ID,32'b10100100011000010001000000000000,MA,32'b11111111111111111111111111111111,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 20
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(20,IA,32'b10000000000000000000000010101000,ID,32'b11010000011000111111111111111111,MA,32'b00000000000000000000000000000001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 21
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(21,IA,32'b10000000000000000000000010101100,ID,32'b01110111111000110000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 22
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(22,IA,32'b10000000000000000000000010111000,ID,32'b10011000011000010001000000000000,MA,32'b00000000000000000000000000000001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 23
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(23,IA,32'b10000000000000000000000010111100,ID,32'b01110111111000110000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 24
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(24,IA,32'b10000000000000000000000011001000,ID,32'b10011000011000100000100000000000,MA,32'b00000000000000000000000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 25
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(25,IA,32'b10000000000000000000000011001100,ID,32'b01110011111000110000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 26
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(26,IA,32'b10000000000000000000000011011000,ID,32'b10000000000111111111100000000000,MA,32'b00000000000000000000000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 27
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(27,IA,32'b10000000000000000000000011011100,ID,32'b01110011111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 28
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(28,IA,32'b10000000000000000000000011101000,ID,32'b11000000000111110000000000000000,MA,32'b00000000000000000000000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 29
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(29,IA,32'b10000000000000000000000011101100,ID,32'b01110011111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 30
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(30,IA,32'b10000000000000000000000011111000,ID,32'b10010000001000001111100000000000,MA,32'b00000000000000000000000000000001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 31
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(31,IA,32'b10000000000000000000000011111100,ID,32'b11010000000000010000000000000001,MA,32'b00000000000000000000000000000001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 32
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(32,IA,32'b10000000000000000000000100000000,ID,32'b01110111111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 33
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(33,IA,32'b10000000000000000000000100001100,ID,32'b11110000010000010000000000000001,MA,32'b00000000000000000000000000000010,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 34
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(34,IA,32'b10000000000000000000000100010000,ID,32'b11010000000000100000000000000010,MA,32'b00000000000000000000000000000001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 35
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(35,IA,32'b10000000000000000000000100010100,ID,32'b01110111111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 36
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(36,IA,32'b10000000000000000000000100100000,ID,32'b10000000011000010001000000000000,MA,32'b00000000000000000000000000000011,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 37
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(37,IA,32'b10000000000000000000000100100100,ID,32'b11010000000000110000000000000011,MA,32'b00000000000000000000000000000001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 38
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(38,IA,32'b10000000000000000000000100101000,ID,32'b01110111111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 39
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(39,IA,32'b10000000000000000000000100110100,ID,32'b11000000100000010000000000000011,MA,32'b00000000000000000000000000000100,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 40
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(40,IA,32'b10000000000000000000000100111000,ID,32'b11010000000001000000000000000100,MA,32'b00000000000000000000000000000001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 41
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(41,IA,32'b10000000000000000000000100111100,ID,32'b01110111111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 42
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(42,IA,32'b10000000000000000000000101001000,ID,32'b11101000101111111111111111111111,MA,32'b11111111111111111111111111111111,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 43
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(43,IA,32'b10000000000000000000000101001100,ID,32'b11101000101001011111111111111010,MA,32'b00000000000000000000000000000101,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 44
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(44,IA,32'b10000000000000000000000101010000,ID,32'b11010000000001010000000000000101,MA,32'b00000000000000000000000000000001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 45
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(45,IA,32'b10000000000000000000000101010100,ID,32'b01110111111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 46
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(46,IA,32'b10000000000000000000000101100000,ID,32'b10100100110001000001000000000000,MA,32'b00000000000000000000000000000110,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 47
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(47,IA,32'b10000000000000000000000101100100,ID,32'b11010000000001100000000000000110,MA,32'b00000000000000000000000000000001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 48
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(48,IA,32'b10000000000000000000000101101000,ID,32'b01110111111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 49
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(49,IA,32'b10000000000000000000000101110100,ID,32'b11000100111111110000000000000001,MA,32'b11111111111111111111111111111111,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 50
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(50,IA,32'b10000000000000000000000101111000,ID,32'b11110100111001110000000000011101,MA,32'b00000000000000000000000000000111,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 51
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(51,IA,32'b10000000000000000000000101111100,ID,32'b11010000000001110000000000000111,MA,32'b00000000000000000000000000000001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 52
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(52,IA,32'b10000000000000000000000110000000,ID,32'b01110111111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 53
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(53,IA,32'b10000000000000000000000110001100,ID,32'b10110001000000010001100000000000,MA,32'b00000000000000000000000000001000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 54
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(54,IA,32'b10000000000000000000000110010000,ID,32'b11010000000010000000000000001000,MA,32'b00000000000000000000000000000001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 55
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(55,IA,32'b10000000000000000000000110010100,ID,32'b01110111111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 56
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(56,IA,32'b10000000000000000000000110100000,ID,32'b10011001001010000100000000000000,MA,32'b00000000000000000000000000000001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 57
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(57,IA,32'b10000000000000000000000110100100,ID,32'b11000101001010011111111111111000,MA,32'b00000000000000000000000000001001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 58
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(58,IA,32'b10000000000000000000000110101000,ID,32'b11010000000010010000000000001001,MA,32'b00000000000000000000000000000001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 59
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(59,IA,32'b10000000000000000000000110101100,ID,32'b01110111111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 60
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(60,IA,32'b10000000000000000000000110111000,ID,32'b10101001010010000001000000000000,MA,32'b00000000000000000000000000001010,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 61
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(61,IA,32'b10000000000000000000000110111100,ID,32'b11010000000010100000000000001010,MA,32'b00000000000000000000000000000001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 62
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(62,IA,32'b10000000000000000000000111000000,ID,32'b01110111111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 63
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(63,IA,32'b10000000000000000000000111001100,ID,32'b11100101011000110000000000001000,MA,32'b00000000000000000000000000001011,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 64
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(64,IA,32'b10000000000000000000000111010000,ID,32'b11010000000010110000000000001011,MA,32'b00000000000000000000000000000001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 65
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(65,IA,32'b10000000000000000000000111010100,ID,32'b01110111111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 66
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(66,IA,32'b10000000000000000000000111100000,ID,32'b10000101100111110000100000000000,MA,32'b11111111111111111111111111111111,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 67
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(67,IA,32'b10000000000000000000000111100100,ID,32'b11110101100011000000000000011101,MA,32'b00000000000000000000000000000111,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 68
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(68,IA,32'b10000000000000000000000111101000,ID,32'b10000001100011000010100000000000,MA,32'b00000000000000000000000000001100,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 69
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(69,IA,32'b10000000000000000000000111101100,ID,32'b11010000000011000000000000001100,MA,32'b00000000000000000000000000000001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 70
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(70,IA,32'b10000000000000000000000111110000,ID,32'b01110111111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 71
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(71,IA,32'b10000000000000000000000111111100,ID,32'b10100101101010000010100000000000,MA,32'b00000000000000000000000000001101,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 72
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(72,IA,32'b10000000000000000000001000000000,ID,32'b11010000000011010000000000001101,MA,32'b00000000000000000000000000000001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 73
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(73,IA,32'b10000000000000000000001000000100,ID,32'b01110111111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 74
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(74,IA,32'b10000000000000000000001000010000,ID,32'b10010101110011000110100000000000,MA,32'b00000000000000000000000000000001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 75
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(75,IA,32'b10000000000000000000001000010100,ID,32'b10000001110011010111000000000000,MA,32'b00000000000000000000000000001110,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 76
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(76,IA,32'b10000000000000000000001000011000,ID,32'b11010000000011100000000000001110,MA,32'b00000000000000000000000000000001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 77
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(77,IA,32'b10000000000000000000001000011100,ID,32'b01110111111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 78
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(78,IA,32'b10000000000000000000001000101000,ID,32'b11110001111000010000000000000100,MA,32'b00000000000000000000000000010000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 79
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(79,IA,32'b10000000000000000000001000101100,ID,32'b10000101111011110000100000000000,MA,32'b00000000000000000000000000001111,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 80
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(80,IA,32'b10000000000000000000001000110000,ID,32'b11010000000011110000000000001111,MA,32'b00000000000000000000000000000001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 81
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(81,IA,32'b10000000000000000000001000110100,ID,32'b01110111111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 82
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(82,IA,32'b10000000000000000000001001000000,ID,32'b10110110000011110001000000000000,MA,32'b00000000000000000000000000000011,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 83
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(83,IA,32'b10000000000000000000001001000100,ID,32'b10000010000100000110100000000000,MA,32'b00000000000000000000000000010000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 84
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(84,IA,32'b10000000000000000000001001001000,ID,32'b11010000000100000000000000010000,MA,32'b00000000000000000000000000000001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 85
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(85,IA,32'b10000000000000000000001001001100,ID,32'b01110111111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 86
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(86,IA,32'b10000000000000000000001001011000,ID,32'b11101110001100001111111111111110,MA,32'b00000000000000000000000000010001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 87
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(87,IA,32'b10000000000000000000001001011100,ID,32'b11010000000100010000000000010001,MA,32'b00000000000000000000000000000001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 88
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(88,IA,32'b10000000000000000000001001100000,ID,32'b01110111111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 89
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(89,IA,32'b10000000000000000000001001101100,ID,32'b10100010010011110001000000000000,MA,32'b00000000000000000000000000000010,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 90
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(90,IA,32'b10000000000000000000001001110000,ID,32'b11100110010100100000000000010000,MA,32'b00000000000000000000000000010010,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 91
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(91,IA,32'b10000000000000000000001001110100,ID,32'b11010000000100100000000000010010,MA,32'b00000000000000000000000000000001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 92
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(92,IA,32'b10000000000000000000001001111000,ID,32'b01110111111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 93
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(93,IA,32'b10000000000000000000001010000100,ID,32'b10111010011011000001000000000000,MA,32'b00000000000000000000000000000011,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 94
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(94,IA,32'b10000000000000000000001010001000,ID,32'b10101110011100001001100000000000,MA,32'b11111111111111111111111111101100,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 95
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(95,IA,32'b10000000000000000000001010001100,ID,32'b11101110011100110000000000000000,MA,32'b00000000000000000000000000010011,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 96
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(96,IA,32'b10000000000000000000001010010000,ID,32'b11010000000100110000000000010011,MA,32'b00000000000000000000000000000001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 97
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(97,IA,32'b10000000000000000000001010010100,ID,32'b01110111111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 98
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(98,IA,32'b10000000000000000000001010100000,ID,32'b11000010100111110000000000011111,MA,32'b00000000000000000000000000011111,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 99
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(99,IA,32'b10000000000000000000001010100100,ID,32'b11100010100101000000000000010100,MA,32'b00000000000000000000000000010100,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 100
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(100,IA,32'b10000000000000000000001010101000,ID,32'b11010000000101000000000000010100,MA,32'b00000000000000000000000000000001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 101
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(101,IA,32'b10000000000000000000001010101100,ID,32'b01110111111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 102
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(102,IA,32'b10000000000000000000001010111000,ID,32'b11100110101101000000000000000001,MA,32'b00000000000000000000000000010101,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 103
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(103,IA,32'b10000000000000000000001010111100,ID,32'b11010000000101010000000000010101,MA,32'b00000000000000000000000000000001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 104
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(104,IA,32'b10000000000000000000001011000000,ID,32'b01110111111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 105
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(105,IA,32'b10000000000000000000001011001100,ID,32'b11000010110100010000000000000101,MA,32'b00000000000000000000000000010110,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 106
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(106,IA,32'b10000000000000000000001011010000,ID,32'b11010000000101100000000000010110,MA,32'b00000000000000000000000000000001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 107
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(107,IA,32'b10000000000000000000001011010100,ID,32'b01110111111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 108
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(108,IA,32'b10000000000000000000001011100000,ID,32'b10101010111101100000100000000000,MA,32'b00000000000000000000000000010111,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 109
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(109,IA,32'b10000000000000000000001011100100,ID,32'b11010000000101110000000000010111,MA,32'b00000000000000000000000000000001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 110
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(110,IA,32'b10000000000000000000001011101000,ID,32'b01110111111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 111
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(111,IA,32'b10000000000000000000001011110100,ID,32'b11100011000101110000000011111100,MA,32'b00000000000000000000000000010100,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 112
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(112,IA,32'b10000000000000000000001011111000,ID,32'b10000011000110000010000000000000,MA,32'b00000000000000000000000000011000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 113
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(113,IA,32'b10000000000000000000001011111100,ID,32'b11010000000110000000000000011000,MA,32'b00000000000000000000000000000001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 114
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(114,IA,32'b10000000000000000000001100000000,ID,32'b01110111111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 115
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(115,IA,32'b10000000000000000000001100001100,ID,32'b10000011001101111100000000000000,MA,32'b00000000000000000000000000101111,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 116
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(116,IA,32'b10000000000000000000001100010000,ID,32'b11000011001110011111111111101010,MA,32'b00000000000000000000000000011001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 117
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(117,IA,32'b10000000000000000000001100010100,ID,32'b11010000000110010000000000011001,MA,32'b00000000000000000000000000000001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 118
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(118,IA,32'b10000000000000000000001100011000,ID,32'b01110111111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 119
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(119,IA,32'b10000000000000000000001100100100,ID,32'b10110011010000110001100000000000,MA,32'b00000000000000000000000000011000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 120
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(120,IA,32'b10000000000000000000001100101000,ID,32'b10100111010000101101000000000000,MA,32'b00000000000000000000000000011010,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 121
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(121,IA,32'b10000000000000000000001100101100,ID,32'b11010000000110100000000000011010,MA,32'b00000000000000000000000000000001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 122
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(122,IA,32'b10000000000000000000001100110000,ID,32'b01110111111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 123
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(123,IA,32'b10000000000000000000001100111100,ID,32'b10000011011011100110100000000000,MA,32'b00000000000000000000000000011011,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 124
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(124,IA,32'b10000000000000000000001101000000,ID,32'b11010000000110110000000000011011,MA,32'b00000000000000000000000000000001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 125
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(125,IA,32'b10000000000000000000001101000100,ID,32'b01110111111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 126
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(126,IA,32'b10000000000000000000001101010000,ID,32'b11000111100101111111111111111011,MA,32'b00000000000000000000000000011100,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 127
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(127,IA,32'b10000000000000000000001101010100,ID,32'b11010000000111000000000000011100,MA,32'b00000000000000000000000000000001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 128
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(128,IA,32'b10000000000000000000001101011000,ID,32'b01110111111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 129
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(129,IA,32'b10000000000000000000001101100100,ID,32'b11000111101111111111111111100011,MA,32'b00000000000000000000000000011101,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 130
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(130,IA,32'b10000000000000000000001101101000,ID,32'b11010000000111010000000000011101,MA,32'b00000000000000000000000000000001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 131
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(131,IA,32'b10000000000000000000001101101100,ID,32'b01110111111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 132
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(132,IA,32'b10000000000000000000001101111000,ID,32'b11000011110111110000000000011111,MA,32'b00000000000000000000000000011111,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 133
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(133,IA,32'b10000000000000000000001101111100,ID,32'b11110111110111100000000000000001,MA,32'b00000000000000000000000000001111,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 134
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(134,IA,32'b10000000000000000000001110000000,ID,32'b11110011110111100000000000000001,MA,32'b00000000000000000000000000011110,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 135
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(135,IA,32'b10000000000000000000001110000100,ID,32'b11010000000111100000000000011110,MA,32'b00000000000000000000000000000001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 136
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(136,IA,32'b10000000000000000000001110001000,ID,32'b01110111111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 137
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(137,IA,32'b10000000000000000000001110010100,ID,32'b01110000000000001111111100011101,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 138
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(138,IA,32'b10000000000000000000001110011000,ID,32'b11000011111111100000000000010001,MA,32'b00000000000000000000000000101111,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 139
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(139,IA,32'b10000000000000000000001110011100,ID,32'b01110011111111110000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 140
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(140,IA,32'b10000000000000000000001110101000,ID,32'b11000010001111110000001111000100,MA,32'b00000000000000000000001111000100,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 141
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(141,IA,32'b10000000000000000000001110101100,ID,32'b11110000001000010000000000011111,MA,32'b10000000000000000000000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 142
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(142,IA,32'b10000000000000000000001110110000,ID,32'b10100110001000011000100000000000,MA,32'b10000000000000000000001111000100,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 143
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(143,IA,32'b10000000000000000000001110110100,ID,32'b01101111100100010000000000000000,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 144
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(144,IA,32'b10000000000000000000001111000100,ID,32'b11110011100111000000000000000001,MA,32'b00000000000000000000011101110000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 145
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(145,IA,32'b10000000000000000000001111001000,ID,32'b11110111100111000000000000000001,MA,32'b00000000000000000000001110111000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 146
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(146,IA,32'b10000000000000000000001111001100,ID,32'b11010010111111000000001110111000,MA,32'b00000000000000000000000000000001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 147
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(147,IA,32'b10000000000000000000001111010000,ID,32'b01110111111101110000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 148
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(148,IA,32'b10000000000000000000001111011100,ID,32'b01111111000111110000000011000000,MA,32'b00000000000000000000011011100000,MOE,1'b1,MWR,1'b0,MRD,32'b10101010101010101010101010101010,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 149
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(149,IA,32'b10000000000000000000001111100000,ID,32'b01111111001111110000000011000000,MA,32'b00000000000000000000011011100100,MOE,1'b1,MWR,1'b0,MRD,32'b01010101010101010101010101010101,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 150
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(150,IA,32'b10000000000000000000001111100100,ID,32'b10000011010110001100100000000000,MA,32'b11111111111111111111111111111111,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 151
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(151,IA,32'b10000000000000000000001111101000,ID,32'b11010011011110101111111111111111,MA,32'b00000000000000000000000000000001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 152
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(152,IA,32'b10000000000000000000001111101100,ID,32'b01110111111110110000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 153
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(153,IA,32'b10000000000000000000001111111000,ID,32'b10000011010110001100000000000000,MA,32'b01010101010101010101010101010100,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 154
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(154,IA,32'b10000000000000000000001111111100,ID,32'b10000111010110101100100000000000,MA,32'b11111111111111111111111111111111,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 155
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(155,IA,32'b10000000000000000000010000000000,ID,32'b11010011011110101111111111111111,MA,32'b00000000000000000000000000000001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 156
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(156,IA,32'b10000000000000000000010000000100,ID,32'b01110111111110110000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 157
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(157,IA,32'b10000000000000000000010000010000,ID,32'b10000011010110011100100000000000,MA,32'b10101010101010101010101010101010,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 158
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(158,IA,32'b10000000000000000000010000010100,ID,32'b10000111010110101100000000000000,MA,32'b00000000000000000000000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 159
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(159,IA,32'b10000000000000000000010000011000,ID,32'b01110011111110100000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 160
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(160,IA,32'b10000000000000000000010000100100,ID,32'b11000010001111110000000000000001,MA,32'b00000000000000000000000000000001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 161
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(161,IA,32'b10000000000000000000010000101000,ID,32'b11000110010100010000000000000001,MA,32'b00000000000000000000000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 162
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(162,IA,32'b10000000000000000000010000101100,ID,32'b01110011111100100000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 163
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(163,IA,32'b10000000000000000000010000111000,ID,32'b11000001011111110000111100001111,MA,32'b00000000000000000000111100001111,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 164
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(164,IA,32'b10000000000000000000010000111100,ID,32'b11000001100111110111111100000000,MA,32'b00000000000000000111111100000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 165
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(165,IA,32'b10000000000000000000010001000000,ID,32'b10100001101010110110000000000000,MA,32'b00000000000000000000111100000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 166
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(166,IA,32'b10000000000000000000010001000100,ID,32'b11010001110011010000111100000000,MA,32'b00000000000000000000000000000001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 167
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(167,IA,32'b10000000000000000000010001001000,ID,32'b01110111111011100000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 168
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(168,IA,32'b10000000000000000000010001010100,ID,32'b10100101101010110110000000000000,MA,32'b00000000000000000111111100001111,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 169
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(169,IA,32'b10000000000000000000010001011000,ID,32'b11010001110011010111111100001111,MA,32'b00000000000000000000000000000001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 170
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(170,IA,32'b10000000000000000000010001011100,ID,32'b01110111111011100000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 171
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(171,IA,32'b10000000000000000000010001101000,ID,32'b10101001101010110110000000000000,MA,32'b00000000000000000111000000001111,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 172
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(172,IA,32'b10000000000000000000010001101100,ID,32'b11010001110011010111000000001111,MA,32'b00000000000000000000000000000001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 173
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(173,IA,32'b10000000000000000000010001110000,ID,32'b01110111111011100000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 174
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(174,IA,32'b10000000000000000000010001111100,ID,32'b10101101101010110110000000000000,MA,32'b11111111111111111000111111110000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 175
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(175,IA,32'b10000000000000000000010010000000,ID,32'b11010001110011011000111111110000,MA,32'b00000000000000000000000000000001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 176
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(176,IA,32'b10000000000000000000010010000100,ID,32'b01110111111011100000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 177
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(177,IA,32'b10000000000000000000010010010000,ID,32'b11000011011111110000000000000001,MA,32'b00000000000000000000000000000001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 178
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(178,IA,32'b10000000000000000000010010010100,ID,32'b11110011100110110000000000100000,MA,32'b00000000000000000000000000000001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 179
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(179,IA,32'b10000000000000000000010010011000,ID,32'b11010011101111000000000000000001,MA,32'b00000000000000000000000000000001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 180
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(180,IA,32'b10000000000000000000010010011100,ID,32'b01110111111111010000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 181
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(181,IA,32'b10000000000000000000010010101000,ID,32'b11110011100110110000000000011111,MA,32'b10000000000000000000000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 182
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(182,IA,32'b10000000000000000000010010101100,ID,32'b11111011010111000000000000010001,MA,32'b11111111111111111100000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 183
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(183,IA,32'b10000000000000000000010010110000,ID,32'b11010011001110101100000000000000,MA,32'b00000000000000000000000000000001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 184
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(184,IA,32'b10000000000000000000010010110100,ID,32'b01110111111110010000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 185
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(185,IA,32'b10000000000000000000010011000000,ID,32'b11110111010111000000000000010001,MA,32'b00000000000000000100000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 186
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(186,IA,32'b10000000000000000000010011000100,ID,32'b11010011001110100100000000000000,MA,32'b00000000000000000000000000000001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 187
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(187,IA,32'b10000000000000000000010011001000,ID,32'b01110111111110010000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 188
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(188,IA,32'b10000000000000000000010011010100,ID,32'b11000011110111110000000000000000,MA,32'b00000000000000000000000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 189
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(189,IA,32'b10000000000000000000010011011000,ID,32'b11000000001111110000000000000000,MA,32'b00000000000000000000000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 190
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(190,IA,32'b10000000000000000000010011011100,ID,32'b00000000000000000000000000010100,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 191
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(191,IA,32'b10000000000000000000000000000100,ID,32'b01110011111111110000000000000011,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 192
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(192,IA,32'b10000000000000000000000000010100,ID,32'b11010000000111100000000000000100,MA,32'b00000000000000000000000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 193
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(193,IA,32'b10000000000000000000000000011000,ID,32'b01110011111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 194
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(194,IA,32'b10000000000000000000000000100100,ID,32'b11000000001000010000000000000001,MA,32'b00000000000000000000000000000001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 195
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(195,IA,32'b10000000000000000000000000101000,ID,32'b01101111111111100000000000000000,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 196
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(196,IA,32'b10000000000000000000010011100000,ID,32'b11110011110111100000000000000001,MA,32'b00000000000000000000100111000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 197
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(197,IA,32'b10000000000000000000010011100100,ID,32'b11110111110111100000000000000001,MA,32'b00000000000000000000010011100000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 198
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(198,IA,32'b10000000000000000000010011101000,ID,32'b11010000000111100000010011100000,MA,32'b00000000000000000000000000000001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 199
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(199,IA,32'b10000000000000000000010011101100,ID,32'b01110111111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 200
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(200,IA,32'b10000000000000000000010011111000,ID,32'b00000100000000000000000000000000,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 201
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(201,IA,32'b10000000000000000000000000000100,ID,32'b01110011111111110000000000000011,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 202
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(202,IA,32'b10000000000000000000000000010100,ID,32'b11010000000111100000000000000100,MA,32'b00000000000000000000000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 203
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(203,IA,32'b10000000000000000000000000011000,ID,32'b01110011111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 204
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(204,IA,32'b10000000000000000000000000100100,ID,32'b11000000001000010000000000000001,MA,32'b00000000000000000000000000000010,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 205
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(205,IA,32'b10000000000000000000000000101000,ID,32'b01101111111111100000000000000000,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 206
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(206,IA,32'b10000000000000000000010011111100,ID,32'b00001000000000000000000000000000,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 207
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(207,IA,32'b10000000000000000000000000000100,ID,32'b01110011111111110000000000000011,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 208
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(208,IA,32'b10000000000000000000000000010100,ID,32'b11010000000111100000000000000100,MA,32'b00000000000000000000000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 209
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(209,IA,32'b10000000000000000000000000011000,ID,32'b01110011111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 210
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(210,IA,32'b10000000000000000000000000100100,ID,32'b11000000001000010000000000000001,MA,32'b00000000000000000000000000000011,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 211
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(211,IA,32'b10000000000000000000000000101000,ID,32'b01101111111111100000000000000000,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 212
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(212,IA,32'b10000000000000000000010100000000,ID,32'b00001100000000000000000000000000,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 213
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(213,IA,32'b10000000000000000000000000000100,ID,32'b01110011111111110000000000000011,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 214
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(214,IA,32'b10000000000000000000000000010100,ID,32'b11010000000111100000000000000100,MA,32'b00000000000000000000000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 215
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(215,IA,32'b10000000000000000000000000011000,ID,32'b01110011111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 216
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(216,IA,32'b10000000000000000000000000100100,ID,32'b11000000001000010000000000000001,MA,32'b00000000000000000000000000000100,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 217
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(217,IA,32'b10000000000000000000000000101000,ID,32'b01101111111111100000000000000000,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 218
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(218,IA,32'b10000000000000000000010100000100,ID,32'b00010000000000000000000000000000,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 219
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(219,IA,32'b10000000000000000000000000000100,ID,32'b01110011111111110000000000000011,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 220
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(220,IA,32'b10000000000000000000000000010100,ID,32'b11010000000111100000000000000100,MA,32'b00000000000000000000000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 221
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(221,IA,32'b10000000000000000000000000011000,ID,32'b01110011111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 222
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(222,IA,32'b10000000000000000000000000100100,ID,32'b11000000001000010000000000000001,MA,32'b00000000000000000000000000000101,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 223
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(223,IA,32'b10000000000000000000000000101000,ID,32'b01101111111111100000000000000000,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 224
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(224,IA,32'b10000000000000000000010100001000,ID,32'b00010100000000000000000000000000,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 225
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(225,IA,32'b10000000000000000000000000000100,ID,32'b01110011111111110000000000000011,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 226
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(226,IA,32'b10000000000000000000000000010100,ID,32'b11010000000111100000000000000100,MA,32'b00000000000000000000000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 227
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(227,IA,32'b10000000000000000000000000011000,ID,32'b01110011111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 228
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(228,IA,32'b10000000000000000000000000100100,ID,32'b11000000001000010000000000000001,MA,32'b00000000000000000000000000000110,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 229
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(229,IA,32'b10000000000000000000000000101000,ID,32'b01101111111111100000000000000000,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 230
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(230,IA,32'b10000000000000000000010100001100,ID,32'b00011000000000000000000000000000,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 231
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(231,IA,32'b10000000000000000000000000000100,ID,32'b01110011111111110000000000000011,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 232
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(232,IA,32'b10000000000000000000000000010100,ID,32'b11010000000111100000000000000100,MA,32'b00000000000000000000000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 233
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(233,IA,32'b10000000000000000000000000011000,ID,32'b01110011111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 234
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(234,IA,32'b10000000000000000000000000100100,ID,32'b11000000001000010000000000000001,MA,32'b00000000000000000000000000000111,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 235
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(235,IA,32'b10000000000000000000000000101000,ID,32'b01101111111111100000000000000000,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 236
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(236,IA,32'b10000000000000000000010100010000,ID,32'b00011100000000000000000000000000,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 237
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(237,IA,32'b10000000000000000000000000000100,ID,32'b01110011111111110000000000000011,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 238
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(238,IA,32'b10000000000000000000000000010100,ID,32'b11010000000111100000000000000100,MA,32'b00000000000000000000000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 239
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(239,IA,32'b10000000000000000000000000011000,ID,32'b01110011111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 240
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(240,IA,32'b10000000000000000000000000100100,ID,32'b11000000001000010000000000000001,MA,32'b00000000000000000000000000001000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 241
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(241,IA,32'b10000000000000000000000000101000,ID,32'b01101111111111100000000000000000,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 242
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(242,IA,32'b10000000000000000000010100010100,ID,32'b00100000000000000000000000000000,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 243
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(243,IA,32'b10000000000000000000000000000100,ID,32'b01110011111111110000000000000011,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 244
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(244,IA,32'b10000000000000000000000000010100,ID,32'b11010000000111100000000000000100,MA,32'b00000000000000000000000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 245
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(245,IA,32'b10000000000000000000000000011000,ID,32'b01110011111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 246
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(246,IA,32'b10000000000000000000000000100100,ID,32'b11000000001000010000000000000001,MA,32'b00000000000000000000000000001001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 247
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(247,IA,32'b10000000000000000000000000101000,ID,32'b01101111111111100000000000000000,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 248
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(248,IA,32'b10000000000000000000010100011000,ID,32'b00100100000000000000000000000000,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 249
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(249,IA,32'b10000000000000000000000000000100,ID,32'b01110011111111110000000000000011,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 250
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(250,IA,32'b10000000000000000000000000010100,ID,32'b11010000000111100000000000000100,MA,32'b00000000000000000000000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 251
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(251,IA,32'b10000000000000000000000000011000,ID,32'b01110011111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 252
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(252,IA,32'b10000000000000000000000000100100,ID,32'b11000000001000010000000000000001,MA,32'b00000000000000000000000000001010,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 253
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(253,IA,32'b10000000000000000000000000101000,ID,32'b01101111111111100000000000000000,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 254
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(254,IA,32'b10000000000000000000010100011100,ID,32'b00101000000000000000000000000000,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 255
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(255,IA,32'b10000000000000000000000000000100,ID,32'b01110011111111110000000000000011,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 256
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(256,IA,32'b10000000000000000000000000010100,ID,32'b11010000000111100000000000000100,MA,32'b00000000000000000000000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 257
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(257,IA,32'b10000000000000000000000000011000,ID,32'b01110011111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 258
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(258,IA,32'b10000000000000000000000000100100,ID,32'b11000000001000010000000000000001,MA,32'b00000000000000000000000000001011,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 259
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(259,IA,32'b10000000000000000000000000101000,ID,32'b01101111111111100000000000000000,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 260
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(260,IA,32'b10000000000000000000010100100000,ID,32'b00101100000000000000000000000000,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 261
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(261,IA,32'b10000000000000000000000000000100,ID,32'b01110011111111110000000000000011,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 262
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(262,IA,32'b10000000000000000000000000010100,ID,32'b11010000000111100000000000000100,MA,32'b00000000000000000000000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 263
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(263,IA,32'b10000000000000000000000000011000,ID,32'b01110011111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 264
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(264,IA,32'b10000000000000000000000000100100,ID,32'b11000000001000010000000000000001,MA,32'b00000000000000000000000000001100,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 265
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(265,IA,32'b10000000000000000000000000101000,ID,32'b01101111111111100000000000000000,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 266
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(266,IA,32'b10000000000000000000010100100100,ID,32'b00110000000000000000000000000000,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 267
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(267,IA,32'b10000000000000000000000000000100,ID,32'b01110011111111110000000000000011,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 268
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(268,IA,32'b10000000000000000000000000010100,ID,32'b11010000000111100000000000000100,MA,32'b00000000000000000000000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 269
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(269,IA,32'b10000000000000000000000000011000,ID,32'b01110011111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 270
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(270,IA,32'b10000000000000000000000000100100,ID,32'b11000000001000010000000000000001,MA,32'b00000000000000000000000000001101,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 271
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(271,IA,32'b10000000000000000000000000101000,ID,32'b01101111111111100000000000000000,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 272
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(272,IA,32'b10000000000000000000010100101000,ID,32'b00110100000000000000000000000000,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 273
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(273,IA,32'b10000000000000000000000000000100,ID,32'b01110011111111110000000000000011,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 274
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(274,IA,32'b10000000000000000000000000010100,ID,32'b11010000000111100000000000000100,MA,32'b00000000000000000000000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 275
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(275,IA,32'b10000000000000000000000000011000,ID,32'b01110011111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 276
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(276,IA,32'b10000000000000000000000000100100,ID,32'b11000000001000010000000000000001,MA,32'b00000000000000000000000000001110,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 277
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(277,IA,32'b10000000000000000000000000101000,ID,32'b01101111111111100000000000000000,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 278
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(278,IA,32'b10000000000000000000010100101100,ID,32'b00111000000000000000000000000000,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 279
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(279,IA,32'b10000000000000000000000000000100,ID,32'b01110011111111110000000000000011,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 280
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(280,IA,32'b10000000000000000000000000010100,ID,32'b11010000000111100000000000000100,MA,32'b00000000000000000000000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 281
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(281,IA,32'b10000000000000000000000000011000,ID,32'b01110011111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 282
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(282,IA,32'b10000000000000000000000000100100,ID,32'b11000000001000010000000000000001,MA,32'b00000000000000000000000000001111,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 283
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(283,IA,32'b10000000000000000000000000101000,ID,32'b01101111111111100000000000000000,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 284
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(284,IA,32'b10000000000000000000010100110000,ID,32'b00111100000000000000000000000000,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 285
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(285,IA,32'b10000000000000000000000000000100,ID,32'b01110011111111110000000000000011,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 286
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(286,IA,32'b10000000000000000000000000010100,ID,32'b11010000000111100000000000000100,MA,32'b00000000000000000000000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 287
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(287,IA,32'b10000000000000000000000000011000,ID,32'b01110011111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 288
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(288,IA,32'b10000000000000000000000000100100,ID,32'b11000000001000010000000000000001,MA,32'b00000000000000000000000000010000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 289
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(289,IA,32'b10000000000000000000000000101000,ID,32'b01101111111111100000000000000000,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 290
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(290,IA,32'b10000000000000000000010100110100,ID,32'b01000000000000000000000000000000,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 291
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(291,IA,32'b10000000000000000000000000000100,ID,32'b01110011111111110000000000000011,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 292
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(292,IA,32'b10000000000000000000000000010100,ID,32'b11010000000111100000000000000100,MA,32'b00000000000000000000000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 293
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(293,IA,32'b10000000000000000000000000011000,ID,32'b01110011111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 294
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(294,IA,32'b10000000000000000000000000100100,ID,32'b11000000001000010000000000000001,MA,32'b00000000000000000000000000010001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 295
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(295,IA,32'b10000000000000000000000000101000,ID,32'b01101111111111100000000000000000,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 296
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(296,IA,32'b10000000000000000000010100111000,ID,32'b01000100000000000000000000000000,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 297
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(297,IA,32'b10000000000000000000000000000100,ID,32'b01110011111111110000000000000011,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 298
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(298,IA,32'b10000000000000000000000000010100,ID,32'b11010000000111100000000000000100,MA,32'b00000000000000000000000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 299
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(299,IA,32'b10000000000000000000000000011000,ID,32'b01110011111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 300
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(300,IA,32'b10000000000000000000000000100100,ID,32'b11000000001000010000000000000001,MA,32'b00000000000000000000000000010010,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 301
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(301,IA,32'b10000000000000000000000000101000,ID,32'b01101111111111100000000000000000,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 302
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(302,IA,32'b10000000000000000000010100111100,ID,32'b01001000000000000000000000000000,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 303
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(303,IA,32'b10000000000000000000000000000100,ID,32'b01110011111111110000000000000011,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 304
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(304,IA,32'b10000000000000000000000000010100,ID,32'b11010000000111100000000000000100,MA,32'b00000000000000000000000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 305
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(305,IA,32'b10000000000000000000000000011000,ID,32'b01110011111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 306
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(306,IA,32'b10000000000000000000000000100100,ID,32'b11000000001000010000000000000001,MA,32'b00000000000000000000000000010011,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 307
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(307,IA,32'b10000000000000000000000000101000,ID,32'b01101111111111100000000000000000,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 308
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(308,IA,32'b10000000000000000000010101000000,ID,32'b01001100000000000000000000000000,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 309
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(309,IA,32'b10000000000000000000000000000100,ID,32'b01110011111111110000000000000011,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 310
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(310,IA,32'b10000000000000000000000000010100,ID,32'b11010000000111100000000000000100,MA,32'b00000000000000000000000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 311
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(311,IA,32'b10000000000000000000000000011000,ID,32'b01110011111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 312
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(312,IA,32'b10000000000000000000000000100100,ID,32'b11000000001000010000000000000001,MA,32'b00000000000000000000000000010100,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 313
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(313,IA,32'b10000000000000000000000000101000,ID,32'b01101111111111100000000000000000,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 314
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(314,IA,32'b10000000000000000000010101000100,ID,32'b01010000000000000000000000000000,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 315
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(315,IA,32'b10000000000000000000000000000100,ID,32'b01110011111111110000000000000011,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 316
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(316,IA,32'b10000000000000000000000000010100,ID,32'b11010000000111100000000000000100,MA,32'b00000000000000000000000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 317
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(317,IA,32'b10000000000000000000000000011000,ID,32'b01110011111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 318
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(318,IA,32'b10000000000000000000000000100100,ID,32'b11000000001000010000000000000001,MA,32'b00000000000000000000000000010101,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 319
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(319,IA,32'b10000000000000000000000000101000,ID,32'b01101111111111100000000000000000,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 320
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(320,IA,32'b10000000000000000000010101001000,ID,32'b01010100000000000000000000000000,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 321
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(321,IA,32'b10000000000000000000000000000100,ID,32'b01110011111111110000000000000011,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 322
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(322,IA,32'b10000000000000000000000000010100,ID,32'b11010000000111100000000000000100,MA,32'b00000000000000000000000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 323
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(323,IA,32'b10000000000000000000000000011000,ID,32'b01110011111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 324
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(324,IA,32'b10000000000000000000000000100100,ID,32'b11000000001000010000000000000001,MA,32'b00000000000000000000000000010110,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 325
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(325,IA,32'b10000000000000000000000000101000,ID,32'b01101111111111100000000000000000,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 326
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(326,IA,32'b10000000000000000000010101001100,ID,32'b01011000000000000000000000000000,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 327
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(327,IA,32'b10000000000000000000000000000100,ID,32'b01110011111111110000000000000011,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 328
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(328,IA,32'b10000000000000000000000000010100,ID,32'b11010000000111100000000000000100,MA,32'b00000000000000000000000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 329
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(329,IA,32'b10000000000000000000000000011000,ID,32'b01110011111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 330
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(330,IA,32'b10000000000000000000000000100100,ID,32'b11000000001000010000000000000001,MA,32'b00000000000000000000000000010111,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 331
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(331,IA,32'b10000000000000000000000000101000,ID,32'b01101111111111100000000000000000,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 332
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(332,IA,32'b10000000000000000000010101010000,ID,32'b01011100000000000000000000000000,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 333
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(333,IA,32'b10000000000000000000000000000100,ID,32'b01110011111111110000000000000011,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 334
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(334,IA,32'b10000000000000000000000000010100,ID,32'b11010000000111100000000000000100,MA,32'b00000000000000000000000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 335
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(335,IA,32'b10000000000000000000000000011000,ID,32'b01110011111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 336
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(336,IA,32'b10000000000000000000000000100100,ID,32'b11000000001000010000000000000001,MA,32'b00000000000000000000000000011000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 337
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(337,IA,32'b10000000000000000000000000101000,ID,32'b01101111111111100000000000000000,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 338
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(338,IA,32'b10000000000000000000010101010100,ID,32'b01101000000000000000000000000000,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 339
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(339,IA,32'b10000000000000000000000000000100,ID,32'b01110011111111110000000000000011,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 340
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(340,IA,32'b10000000000000000000000000010100,ID,32'b11010000000111100000000000000100,MA,32'b00000000000000000000000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 341
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(341,IA,32'b10000000000000000000000000011000,ID,32'b01110011111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 342
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(342,IA,32'b10000000000000000000000000100100,ID,32'b11000000001000010000000000000001,MA,32'b00000000000000000000000000011001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 343
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(343,IA,32'b10000000000000000000000000101000,ID,32'b01101111111111100000000000000000,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 344
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(344,IA,32'b10000000000000000000010101011000,ID,32'b01111000000000000000000000000000,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 345
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(345,IA,32'b10000000000000000000000000000100,ID,32'b01110011111111110000000000000011,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 346
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(346,IA,32'b10000000000000000000000000010100,ID,32'b11010000000111100000000000000100,MA,32'b00000000000000000000000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 347
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(347,IA,32'b10000000000000000000000000011000,ID,32'b01110011111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 348
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(348,IA,32'b10000000000000000000000000100100,ID,32'b11000000001000010000000000000001,MA,32'b00000000000000000000000000011010,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 349
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(349,IA,32'b10000000000000000000000000101000,ID,32'b01101111111111100000000000000000,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 350
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(350,IA,32'b10000000000000000000010101011100,ID,32'b10011100000000000000000000000000,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 351
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(351,IA,32'b10000000000000000000000000000100,ID,32'b01110011111111110000000000000011,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 352
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(352,IA,32'b10000000000000000000000000010100,ID,32'b11010000000111100000000000000100,MA,32'b00000000000000000000000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 353
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(353,IA,32'b10000000000000000000000000011000,ID,32'b01110011111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 354
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(354,IA,32'b10000000000000000000000000100100,ID,32'b11000000001000010000000000000001,MA,32'b00000000000000000000000000011011,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 355
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(355,IA,32'b10000000000000000000000000101000,ID,32'b01101111111111100000000000000000,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 356
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(356,IA,32'b10000000000000000000010101100000,ID,32'b10111100000000000000000000000000,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 357
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(357,IA,32'b10000000000000000000000000000100,ID,32'b01110011111111110000000000000011,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 358
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(358,IA,32'b10000000000000000000000000010100,ID,32'b11010000000111100000000000000100,MA,32'b00000000000000000000000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 359
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(359,IA,32'b10000000000000000000000000011000,ID,32'b01110011111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 360
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(360,IA,32'b10000000000000000000000000100100,ID,32'b11000000001000010000000000000001,MA,32'b00000000000000000000000000011100,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 361
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(361,IA,32'b10000000000000000000000000101000,ID,32'b01101111111111100000000000000000,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 362
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(362,IA,32'b10000000000000000000010101100100,ID,32'b11011100000000000000000000000000,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 363
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(363,IA,32'b10000000000000000000000000000100,ID,32'b01110011111111110000000000000011,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 364
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(364,IA,32'b10000000000000000000000000010100,ID,32'b11010000000111100000000000000100,MA,32'b00000000000000000000000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 365
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(365,IA,32'b10000000000000000000000000011000,ID,32'b01110011111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 366
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(366,IA,32'b10000000000000000000000000100100,ID,32'b11000000001000010000000000000001,MA,32'b00000000000000000000000000011101,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 367
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(367,IA,32'b10000000000000000000000000101000,ID,32'b01101111111111100000000000000000,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 368
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(368,IA,32'b10000000000000000000010101101000,ID,32'b11111100000000000000000000000000,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 369
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(369,IA,32'b10000000000000000000000000000100,ID,32'b01110011111111110000000000000011,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 370
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(370,IA,32'b10000000000000000000000000010100,ID,32'b11010000000111100000000000000100,MA,32'b00000000000000000000000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 371
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(371,IA,32'b10000000000000000000000000011000,ID,32'b01110011111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 372
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(372,IA,32'b10000000000000000000000000100100,ID,32'b11000000001000010000000000000001,MA,32'b00000000000000000000000000011110,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 373
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(373,IA,32'b10000000000000000000000000101000,ID,32'b01101111111111100000000000000000,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 374
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(374,IA,32'b10000000000000000000010101101100,ID,32'b11010000000000010000000000011110,MA,32'b00000000000000000000000000000001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 375
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(375,IA,32'b10000000000000000000010101110000,ID,32'b01110111111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 376
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(376,IA,32'b10000000000000000000010101111100,ID,32'b11000000100111110000011011101000,MA,32'b00000000000000000000011011101000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 377
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(377,IA,32'b10000000000000000000010110000000,ID,32'b01111101001111110000000001010111,MA,32'b00000000000000000000011011100000,MOE,1'b1,MWR,1'b0,MRD,32'b10101010101010101010101010101010,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 378
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(378,IA,32'b10000000000000000000010110000100,ID,32'b11101000000010011111111111111111,MA,32'b01010101010101010101010101010101,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 379
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(379,IA,32'b10000000000000000000010110001000,ID,32'b01100101001001000000000000000000,MA,32'b00000000000000000000011011101000,MOE,1'b0,MWR,1'b1,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'b10101010101010101010101010101010);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 380
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(380,IA,32'b10000000000000000000010110001100,ID,32'b01100100000111110000011011101100,MA,32'b00000000000000000000011011101100,MOE,1'b0,MWR,1'b1,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'b01010101010101010101010101010101);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 381
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(381,IA,32'b10000000000000000000010110010000,ID,32'b01100101001001000000000000001000,MA,32'b00000000000000000000011011110000,MOE,1'b0,MWR,1'b1,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'b10101010101010101010101010101010);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 382
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(382,IA,32'b10000000000000000000010110010100,ID,32'b01100100000111110000011011110100,MA,32'b00000000000000000000011011110100,MOE,1'b0,MWR,1'b1,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'b01010101010101010101010101010101);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 383
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(383,IA,32'b10000000000000000000010110011000,ID,32'b01100000110001000000000000000000,MA,32'b00000000000000000000011011101000,MOE,1'b1,MWR,1'b0,MRD,32'b10101010101010101010101010101010,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 384
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(384,IA,32'b10000000000000000000010110011100,ID,32'b01111100101111110000000001010001,MA,32'b00000000000000000000011011100100,MOE,1'b1,MWR,1'b0,MRD,32'b01010101010101010101010101010101,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 385
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(385,IA,32'b10000000000000000000010110100000,ID,32'b10010000000001100100100000000000,MA,32'b00000000000000000000000000000001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 386
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(386,IA,32'b10000000000000000000010110100100,ID,32'b01110111111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 387
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(387,IA,32'b10000000000000000000010110110000,ID,32'b01100000111111110000011011101100,MA,32'b00000000000000000000011011101100,MOE,1'b1,MWR,1'b0,MRD,32'b01010101010101010101010101010101,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 388
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(388,IA,32'b10000000000000000000010110110100,ID,32'b10010000000001110010100000000000,MA,32'b00000000000000000000000000000001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 389
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(389,IA,32'b10000000000000000000010110111000,ID,32'b01110111111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 390
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(390,IA,32'b10000000000000000000010111000100,ID,32'b01100001000001000000000000001000,MA,32'b00000000000000000000011011110000,MOE,1'b1,MWR,1'b0,MRD,32'b10101010101010101010101010101010,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 391
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(391,IA,32'b10000000000000000000010111001000,ID,32'b10010000000010000100100000000000,MA,32'b00000000000000000000000000000001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 392
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(392,IA,32'b10000000000000000000010111001100,ID,32'b01110111111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 393
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(393,IA,32'b10000000000000000000010111011000,ID,32'b01100001001111110000011011110100,MA,32'b00000000000000000000011011110100,MOE,1'b1,MWR,1'b0,MRD,32'b01010101010101010101010101010101,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 394
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(394,IA,32'b10000000000000000000010111011100,ID,32'b10010000000010010010100000000000,MA,32'b00000000000000000000000000000001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 395
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(395,IA,32'b10000000000000000000010111100000,ID,32'b01110111111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 396
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(396,IA,32'b10000000000000000000010111101100,ID,32'b10000000000111111010000000000000,MA,32'b00000000000000000000000000010100,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 397
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(397,IA,32'b10000000000000000000010111110000,ID,32'b10000000001000000000000000000000,MA,32'b00000000000000000000000000101000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 398
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(398,IA,32'b10000000000000000000010111110100,ID,32'b10000000010000000000000000000000,MA,32'b00000000000000000000000000101000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 399
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(399,IA,32'b10000000000000000000010111111000,ID,32'b10000000011000000000000000000000,MA,32'b00000000000000000000000000101000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 400
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(400,IA,32'b10000000000000000000010111111100,ID,32'b10000000100000000000000000000000,MA,32'b00000000000000000000000000101000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 401
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(401,IA,32'b10000000000000000000011000000000,ID,32'b10000000101000010001000000000000,MA,32'b00000000000000000000000001010000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 402
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(402,IA,32'b10000000000000000000011000000100,ID,32'b10000000101000110010100000000000,MA,32'b00000000000000000000000001111000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 403
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(403,IA,32'b10000000000000000000011000001000,ID,32'b10000000101001000010100000000000,MA,32'b00000000000000000000000010100000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 404
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(404,IA,32'b10000000000000000000011000001100,ID,32'b11010000000001010000000010100000,MA,32'b00000000000000000000000000000001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 405
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(405,IA,32'b10000000000000000000011000010000,ID,32'b01110111111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 406
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(406,IA,32'b10000000000000000000011000011100,ID,32'b01110100000111110000000000000000,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 407
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(407,IA,32'b10000000000000000000011000100000,ID,32'b10000000001000000000000000000000,MA,32'b00000000000000000000110001000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 408
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(408,IA,32'b10000000000000000000011000100100,ID,32'b10000000010000000000000000000000,MA,32'b00000000000000000000110001000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 409
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(409,IA,32'b10000000000000000000011000101000,ID,32'b10000000011000000000000000000000,MA,32'b00000000000000000000110001000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 410
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(410,IA,32'b10000000000000000000011000101100,ID,32'b10000000100000000000000000000000,MA,32'b00000000000000000000110001000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 411
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(411,IA,32'b10000000000000000000011000110000,ID,32'b10000000101000010001000000000000,MA,32'b00000000000000000001100010000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 412
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(412,IA,32'b10000000000000000000011000110100,ID,32'b10000000101000110010100000000000,MA,32'b00000000000000000010010011000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 413
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(413,IA,32'b10000000000000000000011000111000,ID,32'b10000000101001000010100000000000,MA,32'b00000000000000000011000100000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 414
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(414,IA,32'b10000000000000000000011000111100,ID,32'b11010000000001010011000100000000,MA,32'b00000000000000000000000000000001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 415
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(415,IA,32'b10000000000000000000011001000000,ID,32'b01110111111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 416
  RESET=1'b0;
  IRQ=1'b1;
  #1;PRINT(416,IA,32'b10000000000000000000011001001100,ID,32'b11000000000111110000011001010100,MA,32'b00000000000000000000011001010100,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 417
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(417,IA,32'b10000000000000000000011001010000,ID,32'b01101111111000000000000000000000,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 418
  RESET=1'b0;
  IRQ=1'b1;
  #1;PRINT(418,IA,32'b00000000000000000000011001010100,ID,32'b01110011111111110000000000000001,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 419
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(419,IA,32'b10000000000000000000000000001000,ID,32'b01101111111111100000000000000000,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 420
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(420,IA,32'b00000000000000000000011001011000,ID,32'b01110011111111110000000000000011,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 421
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(421,IA,32'b00000000000000000000011001101000,ID,32'b11010000000111100000011001011000,MA,32'b00000000000000000000000000000001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 422
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(422,IA,32'b00000000000000000000011001101100,ID,32'b01110111111000000000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 423
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(423,IA,32'b00000000000000000000011001111000,ID,32'b11000000000111110000011010001100,MA,32'b00000000000000000000011010001100,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 424
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(424,IA,32'b00000000000000000000011001111100,ID,32'b11000000001111110000000000000001,MA,32'b00000000000000000000000000000001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 425
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(425,IA,32'b00000000000000000000011010000000,ID,32'b11110000001000010000000000011111,MA,32'b10000000000000000000000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 426
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(426,IA,32'b00000000000000000000011010000100,ID,32'b10100100000000010000000000000000,MA,32'b10000000000000000000011010001100,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 427
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(427,IA,32'b00000000000000000000011010001000,ID,32'b01101100001000000000000000000000,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 428
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(428,IA,32'b00000000000000000000011010001100,ID,32'b01110000000111110000000000000000,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 429
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(429,IA,32'b00000000000000000000011010010000,ID,32'b11010000001000000000011010010000,MA,32'b00000000000000000000000000000001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 430
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(430,IA,32'b00000000000000000000011010010100,ID,32'b01110111111000010000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 431
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(431,IA,32'b00000000000000000000011010100000,ID,32'b01100000000111110000011011100000,MA,32'b00000000000000000000011011100000,MOE,1'b1,MWR,1'b0,MRD,32'b10101010101010101010101010101010,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 432
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(432,IA,32'b00000000000000000000011010100100,ID,32'b01110011111000000000000000000111,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 433
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(433,IA,32'b00000000000000000000011010101000,ID,32'b01100000000111110000011011100100,MA,32'b00000000000000000000011011100100,MOE,1'b1,MWR,1'b0,MRD,32'b01010101010101010101010101010101,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 434
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(434,IA,32'b00000000000000000000011010101100,ID,32'b01110011111000000000000000000101,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 435
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(435,IA,32'b00000000000000000000011010110000,ID,32'b11000000000111110000000000000000,MA,32'b00000000000000000000000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 436
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(436,IA,32'b00000000000000000000011010110100,ID,32'b01110111111000000000000000000011,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 437
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(437,IA,32'b00000000000000000000011010111000,ID,32'b11000000001111110000000000000001,MA,32'b00000000000000000000000000000001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 438
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(438,IA,32'b00000000000000000000011010111100,ID,32'b11000000010111110000000000100000,MA,32'b00000000000000000000000000100000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 439
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(439,IA,32'b00000000000000000000011011000000,ID,32'b01110111111000010000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 440
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(440,IA,32'b00000000000000000000011011001100,ID,32'b11110000001000010000000000000001,MA,32'b00000000000000000000000000000010,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 441
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(441,IA,32'b00000000000000000000011011010000,ID,32'b11000100010000100000000000000001,MA,32'b00000000000000000000000000011111,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 442
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(442,IA,32'b00000000000000000000011011010100,ID,32'b01110111111000101111111111111010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 443
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(443,IA,32'b00000000000000000000011011000000,ID,32'b01110111111000010000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 444
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(444,IA,32'b00000000000000000000011011001100,ID,32'b11110000001000010000000000000001,MA,32'b00000000000000000000000000000100,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 445
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(445,IA,32'b00000000000000000000011011010000,ID,32'b11000100010000100000000000000001,MA,32'b00000000000000000000000000011110,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 446
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(446,IA,32'b00000000000000000000011011010100,ID,32'b01110111111000101111111111111010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 447
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(447,IA,32'b00000000000000000000011011000000,ID,32'b01110111111000010000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 448
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(448,IA,32'b00000000000000000000011011001100,ID,32'b11110000001000010000000000000001,MA,32'b00000000000000000000000000001000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 449
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(449,IA,32'b00000000000000000000011011010000,ID,32'b11000100010000100000000000000001,MA,32'b00000000000000000000000000011101,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 450
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(450,IA,32'b00000000000000000000011011010100,ID,32'b01110111111000101111111111111010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 451
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(451,IA,32'b00000000000000000000011011000000,ID,32'b01110111111000010000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 452
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(452,IA,32'b00000000000000000000011011001100,ID,32'b11110000001000010000000000000001,MA,32'b00000000000000000000000000010000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 453
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(453,IA,32'b00000000000000000000011011010000,ID,32'b11000100010000100000000000000001,MA,32'b00000000000000000000000000011100,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 454
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(454,IA,32'b00000000000000000000011011010100,ID,32'b01110111111000101111111111111010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 455
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(455,IA,32'b00000000000000000000011011000000,ID,32'b01110111111000010000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 456
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(456,IA,32'b00000000000000000000011011001100,ID,32'b11110000001000010000000000000001,MA,32'b00000000000000000000000000100000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 457
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(457,IA,32'b00000000000000000000011011010000,ID,32'b11000100010000100000000000000001,MA,32'b00000000000000000000000000011011,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 458
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(458,IA,32'b00000000000000000000011011010100,ID,32'b01110111111000101111111111111010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 459
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(459,IA,32'b00000000000000000000011011000000,ID,32'b01110111111000010000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 460
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(460,IA,32'b00000000000000000000011011001100,ID,32'b11110000001000010000000000000001,MA,32'b00000000000000000000000001000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 461
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(461,IA,32'b00000000000000000000011011010000,ID,32'b11000100010000100000000000000001,MA,32'b00000000000000000000000000011010,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 462
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(462,IA,32'b00000000000000000000011011010100,ID,32'b01110111111000101111111111111010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 463
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(463,IA,32'b00000000000000000000011011000000,ID,32'b01110111111000010000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 464
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(464,IA,32'b00000000000000000000011011001100,ID,32'b11110000001000010000000000000001,MA,32'b00000000000000000000000010000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 465
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(465,IA,32'b00000000000000000000011011010000,ID,32'b11000100010000100000000000000001,MA,32'b00000000000000000000000000011001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 466
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(466,IA,32'b00000000000000000000011011010100,ID,32'b01110111111000101111111111111010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 467
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(467,IA,32'b00000000000000000000011011000000,ID,32'b01110111111000010000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 468
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(468,IA,32'b00000000000000000000011011001100,ID,32'b11110000001000010000000000000001,MA,32'b00000000000000000000000100000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 469
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(469,IA,32'b00000000000000000000011011010000,ID,32'b11000100010000100000000000000001,MA,32'b00000000000000000000000000011000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 470
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(470,IA,32'b00000000000000000000011011010100,ID,32'b01110111111000101111111111111010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 471
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(471,IA,32'b00000000000000000000011011000000,ID,32'b01110111111000010000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 472
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(472,IA,32'b00000000000000000000011011001100,ID,32'b11110000001000010000000000000001,MA,32'b00000000000000000000001000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 473
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(473,IA,32'b00000000000000000000011011010000,ID,32'b11000100010000100000000000000001,MA,32'b00000000000000000000000000010111,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 474
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(474,IA,32'b00000000000000000000011011010100,ID,32'b01110111111000101111111111111010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 475
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(475,IA,32'b00000000000000000000011011000000,ID,32'b01110111111000010000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 476
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(476,IA,32'b00000000000000000000011011001100,ID,32'b11110000001000010000000000000001,MA,32'b00000000000000000000010000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 477
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(477,IA,32'b00000000000000000000011011010000,ID,32'b11000100010000100000000000000001,MA,32'b00000000000000000000000000010110,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 478
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(478,IA,32'b00000000000000000000011011010100,ID,32'b01110111111000101111111111111010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 479
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(479,IA,32'b00000000000000000000011011000000,ID,32'b01110111111000010000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 480
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(480,IA,32'b00000000000000000000011011001100,ID,32'b11110000001000010000000000000001,MA,32'b00000000000000000000100000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 481
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(481,IA,32'b00000000000000000000011011010000,ID,32'b11000100010000100000000000000001,MA,32'b00000000000000000000000000010101,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 482
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(482,IA,32'b00000000000000000000011011010100,ID,32'b01110111111000101111111111111010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 483
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(483,IA,32'b00000000000000000000011011000000,ID,32'b01110111111000010000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 484
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(484,IA,32'b00000000000000000000011011001100,ID,32'b11110000001000010000000000000001,MA,32'b00000000000000000001000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 485
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(485,IA,32'b00000000000000000000011011010000,ID,32'b11000100010000100000000000000001,MA,32'b00000000000000000000000000010100,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 486
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(486,IA,32'b00000000000000000000011011010100,ID,32'b01110111111000101111111111111010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 487
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(487,IA,32'b00000000000000000000011011000000,ID,32'b01110111111000010000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 488
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(488,IA,32'b00000000000000000000011011001100,ID,32'b11110000001000010000000000000001,MA,32'b00000000000000000010000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 489
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(489,IA,32'b00000000000000000000011011010000,ID,32'b11000100010000100000000000000001,MA,32'b00000000000000000000000000010011,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 490
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(490,IA,32'b00000000000000000000011011010100,ID,32'b01110111111000101111111111111010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 491
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(491,IA,32'b00000000000000000000011011000000,ID,32'b01110111111000010000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 492
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(492,IA,32'b00000000000000000000011011001100,ID,32'b11110000001000010000000000000001,MA,32'b00000000000000000100000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 493
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(493,IA,32'b00000000000000000000011011010000,ID,32'b11000100010000100000000000000001,MA,32'b00000000000000000000000000010010,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 494
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(494,IA,32'b00000000000000000000011011010100,ID,32'b01110111111000101111111111111010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 495
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(495,IA,32'b00000000000000000000011011000000,ID,32'b01110111111000010000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 496
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(496,IA,32'b00000000000000000000011011001100,ID,32'b11110000001000010000000000000001,MA,32'b00000000000000001000000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 497
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(497,IA,32'b00000000000000000000011011010000,ID,32'b11000100010000100000000000000001,MA,32'b00000000000000000000000000010001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 498
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(498,IA,32'b00000000000000000000011011010100,ID,32'b01110111111000101111111111111010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 499
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(499,IA,32'b00000000000000000000011011000000,ID,32'b01110111111000010000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 500
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(500,IA,32'b00000000000000000000011011001100,ID,32'b11110000001000010000000000000001,MA,32'b00000000000000010000000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 501
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(501,IA,32'b00000000000000000000011011010000,ID,32'b11000100010000100000000000000001,MA,32'b00000000000000000000000000010000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 502
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(502,IA,32'b00000000000000000000011011010100,ID,32'b01110111111000101111111111111010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 503
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(503,IA,32'b00000000000000000000011011000000,ID,32'b01110111111000010000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 504
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(504,IA,32'b00000000000000000000011011001100,ID,32'b11110000001000010000000000000001,MA,32'b00000000000000100000000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 505
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(505,IA,32'b00000000000000000000011011010000,ID,32'b11000100010000100000000000000001,MA,32'b00000000000000000000000000001111,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 506
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(506,IA,32'b00000000000000000000011011010100,ID,32'b01110111111000101111111111111010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 507
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(507,IA,32'b00000000000000000000011011000000,ID,32'b01110111111000010000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 508
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(508,IA,32'b00000000000000000000011011001100,ID,32'b11110000001000010000000000000001,MA,32'b00000000000001000000000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 509
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(509,IA,32'b00000000000000000000011011010000,ID,32'b11000100010000100000000000000001,MA,32'b00000000000000000000000000001110,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 510
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(510,IA,32'b00000000000000000000011011010100,ID,32'b01110111111000101111111111111010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 511
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(511,IA,32'b00000000000000000000011011000000,ID,32'b01110111111000010000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 512
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(512,IA,32'b00000000000000000000011011001100,ID,32'b11110000001000010000000000000001,MA,32'b00000000000010000000000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 513
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(513,IA,32'b00000000000000000000011011010000,ID,32'b11000100010000100000000000000001,MA,32'b00000000000000000000000000001101,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 514
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(514,IA,32'b00000000000000000000011011010100,ID,32'b01110111111000101111111111111010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 515
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(515,IA,32'b00000000000000000000011011000000,ID,32'b01110111111000010000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 516
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(516,IA,32'b00000000000000000000011011001100,ID,32'b11110000001000010000000000000001,MA,32'b00000000000100000000000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 517
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(517,IA,32'b00000000000000000000011011010000,ID,32'b11000100010000100000000000000001,MA,32'b00000000000000000000000000001100,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 518
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(518,IA,32'b00000000000000000000011011010100,ID,32'b01110111111000101111111111111010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 519
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(519,IA,32'b00000000000000000000011011000000,ID,32'b01110111111000010000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 520
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(520,IA,32'b00000000000000000000011011001100,ID,32'b11110000001000010000000000000001,MA,32'b00000000001000000000000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 521
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(521,IA,32'b00000000000000000000011011010000,ID,32'b11000100010000100000000000000001,MA,32'b00000000000000000000000000001011,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 522
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(522,IA,32'b00000000000000000000011011010100,ID,32'b01110111111000101111111111111010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 523
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(523,IA,32'b00000000000000000000011011000000,ID,32'b01110111111000010000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 524
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(524,IA,32'b00000000000000000000011011001100,ID,32'b11110000001000010000000000000001,MA,32'b00000000010000000000000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 525
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(525,IA,32'b00000000000000000000011011010000,ID,32'b11000100010000100000000000000001,MA,32'b00000000000000000000000000001010,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 526
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(526,IA,32'b00000000000000000000011011010100,ID,32'b01110111111000101111111111111010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 527
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(527,IA,32'b00000000000000000000011011000000,ID,32'b01110111111000010000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 528
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(528,IA,32'b00000000000000000000011011001100,ID,32'b11110000001000010000000000000001,MA,32'b00000000100000000000000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 529
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(529,IA,32'b00000000000000000000011011010000,ID,32'b11000100010000100000000000000001,MA,32'b00000000000000000000000000001001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 530
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(530,IA,32'b00000000000000000000011011010100,ID,32'b01110111111000101111111111111010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 531
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(531,IA,32'b00000000000000000000011011000000,ID,32'b01110111111000010000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 532
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(532,IA,32'b00000000000000000000011011001100,ID,32'b11110000001000010000000000000001,MA,32'b00000001000000000000000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 533
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(533,IA,32'b00000000000000000000011011010000,ID,32'b11000100010000100000000000000001,MA,32'b00000000000000000000000000001000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 534
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(534,IA,32'b00000000000000000000011011010100,ID,32'b01110111111000101111111111111010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 535
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(535,IA,32'b00000000000000000000011011000000,ID,32'b01110111111000010000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 536
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(536,IA,32'b00000000000000000000011011001100,ID,32'b11110000001000010000000000000001,MA,32'b00000010000000000000000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 537
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(537,IA,32'b00000000000000000000011011010000,ID,32'b11000100010000100000000000000001,MA,32'b00000000000000000000000000000111,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 538
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(538,IA,32'b00000000000000000000011011010100,ID,32'b01110111111000101111111111111010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 539
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(539,IA,32'b00000000000000000000011011000000,ID,32'b01110111111000010000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 540
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(540,IA,32'b00000000000000000000011011001100,ID,32'b11110000001000010000000000000001,MA,32'b00000100000000000000000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 541
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(541,IA,32'b00000000000000000000011011010000,ID,32'b11000100010000100000000000000001,MA,32'b00000000000000000000000000000110,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 542
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(542,IA,32'b00000000000000000000011011010100,ID,32'b01110111111000101111111111111010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 543
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(543,IA,32'b00000000000000000000011011000000,ID,32'b01110111111000010000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 544
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(544,IA,32'b00000000000000000000011011001100,ID,32'b11110000001000010000000000000001,MA,32'b00001000000000000000000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 545
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(545,IA,32'b00000000000000000000011011010000,ID,32'b11000100010000100000000000000001,MA,32'b00000000000000000000000000000101,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 546
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(546,IA,32'b00000000000000000000011011010100,ID,32'b01110111111000101111111111111010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 547
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(547,IA,32'b00000000000000000000011011000000,ID,32'b01110111111000010000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 548
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(548,IA,32'b00000000000000000000011011001100,ID,32'b11110000001000010000000000000001,MA,32'b00010000000000000000000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 549
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(549,IA,32'b00000000000000000000011011010000,ID,32'b11000100010000100000000000000001,MA,32'b00000000000000000000000000000100,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 550
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(550,IA,32'b00000000000000000000011011010100,ID,32'b01110111111000101111111111111010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 551
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(551,IA,32'b00000000000000000000011011000000,ID,32'b01110111111000010000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 552
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(552,IA,32'b00000000000000000000011011001100,ID,32'b11110000001000010000000000000001,MA,32'b00100000000000000000000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 553
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(553,IA,32'b00000000000000000000011011010000,ID,32'b11000100010000100000000000000001,MA,32'b00000000000000000000000000000011,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 554
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(554,IA,32'b00000000000000000000011011010100,ID,32'b01110111111000101111111111111010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 555
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(555,IA,32'b00000000000000000000011011000000,ID,32'b01110111111000010000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 556
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(556,IA,32'b00000000000000000000011011001100,ID,32'b11110000001000010000000000000001,MA,32'b01000000000000000000000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 557
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(557,IA,32'b00000000000000000000011011010000,ID,32'b11000100010000100000000000000001,MA,32'b00000000000000000000000000000010,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 558
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(558,IA,32'b00000000000000000000011011010100,ID,32'b01110111111000101111111111111010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 559
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(559,IA,32'b00000000000000000000011011000000,ID,32'b01110111111000010000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 560
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(560,IA,32'b00000000000000000000011011001100,ID,32'b11110000001000010000000000000001,MA,32'b10000000000000000000000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 561
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(561,IA,32'b00000000000000000000011011010000,ID,32'b11000100010000100000000000000001,MA,32'b00000000000000000000000000000001,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 562
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(562,IA,32'b00000000000000000000011011010100,ID,32'b01110111111000101111111111111010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 563
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(563,IA,32'b00000000000000000000011011000000,ID,32'b01110111111000010000000000000010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 564
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(564,IA,32'b00000000000000000000011011001100,ID,32'b11110000001000010000000000000001,MA,32'b00000000000000000000000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 565
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(565,IA,32'b00000000000000000000011011010000,ID,32'b11000100010000100000000000000001,MA,32'b00000000000000000000000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 566
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(566,IA,32'b00000000000000000000011011010100,ID,32'b01110111111000101111111111111010,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 567
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(567,IA,32'b00000000000000000000011011011000,ID,32'b11000011111111110000000000000000,MA,32'b00000000000000000000000000000000,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;

  //CASE: 568
  RESET=1'b0;
  IRQ=1'b0;
  #1;PRINT(568,IA,32'b00000000000000000000011011011100,ID,32'b01110011111111111111111111111110,MA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MOE,1'bx,MWR,1'b0,MRD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,MWD,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  CLK=1;
  #10;
  CLK=0;


  if(weAreOk) $display("TEST OK\n\nPassed");


  end

endmodule