`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Abdelrahman Elbehery
//
// Create Date:   00:36:55 02/10/2017
// Design Name:   SHIFT
// Module Name:   F:/Self learning/FPGA/Projects/BETA_ISE/TB_SHIFT.v
// Project Name:  BETA_ISE
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: SHIFT
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module TB_SHIFT;
  reg CLK=0;
  integer weAreOk=1;

  task PRINT;
    input integer CN;
    input [31:0] Y;
    input [31:0] ExY;
    if( Y!=ExY ) begin
    $display("Error in case: %d\nY: %b\nExpected: %b\n",CN,Y,ExY);
    weAreOk=0;
    end
  endtask

  reg [1:0] SFN;
  reg [31:0] A;
  reg [4:0] B;
  wire [31:0] Y;

  SHIFT uut(.SFN(SFN),.A(A),.B(B),.Y(Y));



initial begin
  //CASE: 1
  SFN=2'b00;
  A=32'b00000000000000000000000000000000;
  B=5'b00000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(1,Y,32'b00000000000000000000000000000000);
  #10;

  //CASE: 2
  SFN=2'b01;
  A=32'b00000000000000000000000000000000;
  B=5'b00000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(2,Y,32'b00000000000000000000000000000000);
  #10;

  //CASE: 3
  SFN=2'b11;
  A=32'b00000000000000000000000000000000;
  B=5'b00000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(3,Y,32'b00000000000000000000000000000000);
  #10;

  //CASE: 4
  SFN=2'b00;
  A=32'b00000000000000000000000000000000;
  B=5'b00001;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(4,Y,32'b00000000000000000000000000000000);
  #10;

  //CASE: 5
  SFN=2'b01;
  A=32'b00000000000000000000000000000000;
  B=5'b00001;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(5,Y,32'b00000000000000000000000000000000);
  #10;

  //CASE: 6
  SFN=2'b11;
  A=32'b00000000000000000000000000000000;
  B=5'b00001;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(6,Y,32'b00000000000000000000000000000000);
  #10;

  //CASE: 7
  SFN=2'b00;
  A=32'b00000000000000000000000000000000;
  B=5'b00010;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(7,Y,32'b00000000000000000000000000000000);
  #10;

  //CASE: 8
  SFN=2'b01;
  A=32'b00000000000000000000000000000000;
  B=5'b00010;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(8,Y,32'b00000000000000000000000000000000);
  #10;

  //CASE: 9
  SFN=2'b11;
  A=32'b00000000000000000000000000000000;
  B=5'b00010;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(9,Y,32'b00000000000000000000000000000000);
  #10;

  //CASE: 10
  SFN=2'b00;
  A=32'b00000000000000000000000000000000;
  B=5'b00100;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(10,Y,32'b00000000000000000000000000000000);
  #10;

  //CASE: 11
  SFN=2'b01;
  A=32'b00000000000000000000000000000000;
  B=5'b00100;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(11,Y,32'b00000000000000000000000000000000);
  #10;

  //CASE: 12
  SFN=2'b11;
  A=32'b00000000000000000000000000000000;
  B=5'b00100;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(12,Y,32'b00000000000000000000000000000000);
  #10;

  //CASE: 13
  SFN=2'b00;
  A=32'b00000000000000000000000000000000;
  B=5'b01000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(13,Y,32'b00000000000000000000000000000000);
  #10;

  //CASE: 14
  SFN=2'b01;
  A=32'b00000000000000000000000000000000;
  B=5'b01000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(14,Y,32'b00000000000000000000000000000000);
  #10;

  //CASE: 15
  SFN=2'b11;
  A=32'b00000000000000000000000000000000;
  B=5'b01000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(15,Y,32'b00000000000000000000000000000000);
  #10;

  //CASE: 16
  SFN=2'b00;
  A=32'b00000000000000000000000000000000;
  B=5'b10000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(16,Y,32'b00000000000000000000000000000000);
  #10;

  //CASE: 17
  SFN=2'b01;
  A=32'b00000000000000000000000000000000;
  B=5'b10000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(17,Y,32'b00000000000000000000000000000000);
  #10;

  //CASE: 18
  SFN=2'b11;
  A=32'b00000000000000000000000000000000;
  B=5'b10000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(18,Y,32'b00000000000000000000000000000000);
  #10;

  //CASE: 19
  SFN=2'b00;
  A=32'b00000000000000000000000000000000;
  B=5'b11111;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(19,Y,32'b00000000000000000000000000000000);
  #10;

  //CASE: 20
  SFN=2'b01;
  A=32'b00000000000000000000000000000000;
  B=5'b11111;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(20,Y,32'b00000000000000000000000000000000);
  #10;

  //CASE: 21
  SFN=2'b11;
  A=32'b00000000000000000000000000000000;
  B=5'b11111;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(21,Y,32'b00000000000000000000000000000000);
  #10;

  //CASE: 22
  SFN=2'b00;
  A=32'b00000000000000000000000000000001;
  B=5'b00000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(22,Y,32'b00000000000000000000000000000001);
  #10;

  //CASE: 23
  SFN=2'b01;
  A=32'b00000000000000000000000000000001;
  B=5'b00000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(23,Y,32'b00000000000000000000000000000001);
  #10;

  //CASE: 24
  SFN=2'b11;
  A=32'b00000000000000000000000000000001;
  B=5'b00000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(24,Y,32'b00000000000000000000000000000001);
  #10;

  //CASE: 25
  SFN=2'b00;
  A=32'b00000000000000000000000000000001;
  B=5'b00001;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(25,Y,32'b00000000000000000000000000000010);
  #10;

  //CASE: 26
  SFN=2'b01;
  A=32'b00000000000000000000000000000001;
  B=5'b00001;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(26,Y,32'b00000000000000000000000000000000);
  #10;

  //CASE: 27
  SFN=2'b11;
  A=32'b00000000000000000000000000000001;
  B=5'b00001;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(27,Y,32'b00000000000000000000000000000000);
  #10;

  //CASE: 28
  SFN=2'b00;
  A=32'b00000000000000000000000000000001;
  B=5'b00010;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(28,Y,32'b00000000000000000000000000000100);
  #10;

  //CASE: 29
  SFN=2'b01;
  A=32'b00000000000000000000000000000001;
  B=5'b00010;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(29,Y,32'b00000000000000000000000000000000);
  #10;

  //CASE: 30
  SFN=2'b11;
  A=32'b00000000000000000000000000000001;
  B=5'b00010;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(30,Y,32'b00000000000000000000000000000000);
  #10;

  //CASE: 31
  SFN=2'b00;
  A=32'b00000000000000000000000000000001;
  B=5'b00100;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(31,Y,32'b00000000000000000000000000010000);
  #10;

  //CASE: 32
  SFN=2'b01;
  A=32'b00000000000000000000000000000001;
  B=5'b00100;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(32,Y,32'b00000000000000000000000000000000);
  #10;

  //CASE: 33
  SFN=2'b11;
  A=32'b00000000000000000000000000000001;
  B=5'b00100;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(33,Y,32'b00000000000000000000000000000000);
  #10;

  //CASE: 34
  SFN=2'b00;
  A=32'b00000000000000000000000000000001;
  B=5'b01000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(34,Y,32'b00000000000000000000000100000000);
  #10;

  //CASE: 35
  SFN=2'b01;
  A=32'b00000000000000000000000000000001;
  B=5'b01000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(35,Y,32'b00000000000000000000000000000000);
  #10;

  //CASE: 36
  SFN=2'b11;
  A=32'b00000000000000000000000000000001;
  B=5'b01000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(36,Y,32'b00000000000000000000000000000000);
  #10;

  //CASE: 37
  SFN=2'b00;
  A=32'b00000000000000000000000000000001;
  B=5'b10000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(37,Y,32'b00000000000000010000000000000000);
  #10;

  //CASE: 38
  SFN=2'b01;
  A=32'b00000000000000000000000000000001;
  B=5'b10000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(38,Y,32'b00000000000000000000000000000000);
  #10;

  //CASE: 39
  SFN=2'b11;
  A=32'b00000000000000000000000000000001;
  B=5'b10000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(39,Y,32'b00000000000000000000000000000000);
  #10;

  //CASE: 40
  SFN=2'b00;
  A=32'b00000000000000000000000000000001;
  B=5'b11111;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(40,Y,32'b10000000000000000000000000000000);
  #10;

  //CASE: 41
  SFN=2'b01;
  A=32'b00000000000000000000000000000001;
  B=5'b11111;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(41,Y,32'b00000000000000000000000000000000);
  #10;

  //CASE: 42
  SFN=2'b11;
  A=32'b00000000000000000000000000000001;
  B=5'b11111;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(42,Y,32'b00000000000000000000000000000000);
  #10;

  //CASE: 43
  SFN=2'b00;
  A=32'b11111111111111111111111111111111;
  B=5'b00000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(43,Y,32'b11111111111111111111111111111111);
  #10;

  //CASE: 44
  SFN=2'b01;
  A=32'b11111111111111111111111111111111;
  B=5'b00000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(44,Y,32'b11111111111111111111111111111111);
  #10;

  //CASE: 45
  SFN=2'b11;
  A=32'b11111111111111111111111111111111;
  B=5'b00000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(45,Y,32'b11111111111111111111111111111111);
  #10;

  //CASE: 46
  SFN=2'b00;
  A=32'b11111111111111111111111111111111;
  B=5'b00001;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(46,Y,32'b11111111111111111111111111111110);
  #10;

  //CASE: 47
  SFN=2'b01;
  A=32'b11111111111111111111111111111111;
  B=5'b00001;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(47,Y,32'b01111111111111111111111111111111);
  #10;

  //CASE: 48
  SFN=2'b11;
  A=32'b11111111111111111111111111111111;
  B=5'b00001;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(48,Y,32'b11111111111111111111111111111111);
  #10;

  //CASE: 49
  SFN=2'b00;
  A=32'b11111111111111111111111111111111;
  B=5'b00010;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(49,Y,32'b11111111111111111111111111111100);
  #10;

  //CASE: 50
  SFN=2'b01;
  A=32'b11111111111111111111111111111111;
  B=5'b00010;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(50,Y,32'b00111111111111111111111111111111);
  #10;

  //CASE: 51
  SFN=2'b11;
  A=32'b11111111111111111111111111111111;
  B=5'b00010;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(51,Y,32'b11111111111111111111111111111111);
  #10;

  //CASE: 52
  SFN=2'b00;
  A=32'b11111111111111111111111111111111;
  B=5'b00100;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(52,Y,32'b11111111111111111111111111110000);
  #10;

  //CASE: 53
  SFN=2'b01;
  A=32'b11111111111111111111111111111111;
  B=5'b00100;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(53,Y,32'b00001111111111111111111111111111);
  #10;

  //CASE: 54
  SFN=2'b11;
  A=32'b11111111111111111111111111111111;
  B=5'b00100;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(54,Y,32'b11111111111111111111111111111111);
  #10;

  //CASE: 55
  SFN=2'b00;
  A=32'b11111111111111111111111111111111;
  B=5'b01000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(55,Y,32'b11111111111111111111111100000000);
  #10;

  //CASE: 56
  SFN=2'b01;
  A=32'b11111111111111111111111111111111;
  B=5'b01000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(56,Y,32'b00000000111111111111111111111111);
  #10;

  //CASE: 57
  SFN=2'b11;
  A=32'b11111111111111111111111111111111;
  B=5'b01000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(57,Y,32'b11111111111111111111111111111111);
  #10;

  //CASE: 58
  SFN=2'b00;
  A=32'b11111111111111111111111111111111;
  B=5'b10000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(58,Y,32'b11111111111111110000000000000000);
  #10;

  //CASE: 59
  SFN=2'b01;
  A=32'b11111111111111111111111111111111;
  B=5'b10000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(59,Y,32'b00000000000000001111111111111111);
  #10;

  //CASE: 60
  SFN=2'b11;
  A=32'b11111111111111111111111111111111;
  B=5'b10000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(60,Y,32'b11111111111111111111111111111111);
  #10;

  //CASE: 61
  SFN=2'b00;
  A=32'b11111111111111111111111111111111;
  B=5'b11111;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(61,Y,32'b10000000000000000000000000000000);
  #10;

  //CASE: 62
  SFN=2'b01;
  A=32'b11111111111111111111111111111111;
  B=5'b11111;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(62,Y,32'b00000000000000000000000000000001);
  #10;

  //CASE: 63
  SFN=2'b11;
  A=32'b11111111111111111111111111111111;
  B=5'b11111;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(63,Y,32'b11111111111111111111111111111111);
  #10;

  //CASE: 64
  SFN=2'b00;
  A=32'b00010010001101000101011001111000;
  B=5'b00000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(64,Y,32'b00010010001101000101011001111000);
  #10;

  //CASE: 65
  SFN=2'b01;
  A=32'b00010010001101000101011001111000;
  B=5'b00000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(65,Y,32'b00010010001101000101011001111000);
  #10;

  //CASE: 66
  SFN=2'b11;
  A=32'b00010010001101000101011001111000;
  B=5'b00000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(66,Y,32'b00010010001101000101011001111000);
  #10;

  //CASE: 67
  SFN=2'b00;
  A=32'b00010010001101000101011001111000;
  B=5'b00001;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(67,Y,32'b00100100011010001010110011110000);
  #10;

  //CASE: 68
  SFN=2'b01;
  A=32'b00010010001101000101011001111000;
  B=5'b00001;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(68,Y,32'b00001001000110100010101100111100);
  #10;

  //CASE: 69
  SFN=2'b11;
  A=32'b00010010001101000101011001111000;
  B=5'b00001;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(69,Y,32'b00001001000110100010101100111100);
  #10;

  //CASE: 70
  SFN=2'b00;
  A=32'b00010010001101000101011001111000;
  B=5'b00010;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(70,Y,32'b01001000110100010101100111100000);
  #10;

  //CASE: 71
  SFN=2'b01;
  A=32'b00010010001101000101011001111000;
  B=5'b00010;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(71,Y,32'b00000100100011010001010110011110);
  #10;

  //CASE: 72
  SFN=2'b11;
  A=32'b00010010001101000101011001111000;
  B=5'b00010;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(72,Y,32'b00000100100011010001010110011110);
  #10;

  //CASE: 73
  SFN=2'b00;
  A=32'b00010010001101000101011001111000;
  B=5'b00100;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(73,Y,32'b00100011010001010110011110000000);
  #10;

  //CASE: 74
  SFN=2'b01;
  A=32'b00010010001101000101011001111000;
  B=5'b00100;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(74,Y,32'b00000001001000110100010101100111);
  #10;

  //CASE: 75
  SFN=2'b11;
  A=32'b00010010001101000101011001111000;
  B=5'b00100;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(75,Y,32'b00000001001000110100010101100111);
  #10;

  //CASE: 76
  SFN=2'b00;
  A=32'b00010010001101000101011001111000;
  B=5'b01000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(76,Y,32'b00110100010101100111100000000000);
  #10;

  //CASE: 77
  SFN=2'b01;
  A=32'b00010010001101000101011001111000;
  B=5'b01000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(77,Y,32'b00000000000100100011010001010110);
  #10;

  //CASE: 78
  SFN=2'b11;
  A=32'b00010010001101000101011001111000;
  B=5'b01000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(78,Y,32'b00000000000100100011010001010110);
  #10;

  //CASE: 79
  SFN=2'b00;
  A=32'b00010010001101000101011001111000;
  B=5'b10000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(79,Y,32'b01010110011110000000000000000000);
  #10;

  //CASE: 80
  SFN=2'b01;
  A=32'b00010010001101000101011001111000;
  B=5'b10000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(80,Y,32'b00000000000000000001001000110100);
  #10;

  //CASE: 81
  SFN=2'b11;
  A=32'b00010010001101000101011001111000;
  B=5'b10000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(81,Y,32'b00000000000000000001001000110100);
  #10;

  //CASE: 82
  SFN=2'b00;
  A=32'b00010010001101000101011001111000;
  B=5'b11111;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(82,Y,32'b00000000000000000000000000000000);
  #10;

  //CASE: 83
  SFN=2'b01;
  A=32'b00010010001101000101011001111000;
  B=5'b11111;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(83,Y,32'b00000000000000000000000000000000);
  #10;

  //CASE: 84
  SFN=2'b11;
  A=32'b00010010001101000101011001111000;
  B=5'b11111;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(84,Y,32'b00000000000000000000000000000000);
  #10;

  //CASE: 85
  SFN=2'b00;
  A=32'b11111110110111001011101010011000;
  B=5'b00000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(85,Y,32'b11111110110111001011101010011000);
  #10;

  //CASE: 86
  SFN=2'b01;
  A=32'b11111110110111001011101010011000;
  B=5'b00000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(86,Y,32'b11111110110111001011101010011000);
  #10;

  //CASE: 87
  SFN=2'b11;
  A=32'b11111110110111001011101010011000;
  B=5'b00000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(87,Y,32'b11111110110111001011101010011000);
  #10;

  //CASE: 88
  SFN=2'b00;
  A=32'b11111110110111001011101010011000;
  B=5'b00001;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(88,Y,32'b11111101101110010111010100110000);
  #10;

  //CASE: 89
  SFN=2'b01;
  A=32'b11111110110111001011101010011000;
  B=5'b00001;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(89,Y,32'b01111111011011100101110101001100);
  #10;

  //CASE: 90
  SFN=2'b11;
  A=32'b11111110110111001011101010011000;
  B=5'b00001;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(90,Y,32'b11111111011011100101110101001100);
  #10;

  //CASE: 91
  SFN=2'b00;
  A=32'b11111110110111001011101010011000;
  B=5'b00010;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(91,Y,32'b11111011011100101110101001100000);
  #10;

  //CASE: 92
  SFN=2'b01;
  A=32'b11111110110111001011101010011000;
  B=5'b00010;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(92,Y,32'b00111111101101110010111010100110);
  #10;

  //CASE: 93
  SFN=2'b11;
  A=32'b11111110110111001011101010011000;
  B=5'b00010;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(93,Y,32'b11111111101101110010111010100110);
  #10;

  //CASE: 94
  SFN=2'b00;
  A=32'b11111110110111001011101010011000;
  B=5'b00100;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(94,Y,32'b11101101110010111010100110000000);
  #10;

  //CASE: 95
  SFN=2'b01;
  A=32'b11111110110111001011101010011000;
  B=5'b00100;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(95,Y,32'b00001111111011011100101110101001);
  #10;

  //CASE: 96
  SFN=2'b11;
  A=32'b11111110110111001011101010011000;
  B=5'b00100;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(96,Y,32'b11111111111011011100101110101001);
  #10;

  //CASE: 97
  SFN=2'b00;
  A=32'b11111110110111001011101010011000;
  B=5'b01000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(97,Y,32'b11011100101110101001100000000000);
  #10;

  //CASE: 98
  SFN=2'b01;
  A=32'b11111110110111001011101010011000;
  B=5'b01000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(98,Y,32'b00000000111111101101110010111010);
  #10;

  //CASE: 99
  SFN=2'b11;
  A=32'b11111110110111001011101010011000;
  B=5'b01000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(99,Y,32'b11111111111111101101110010111010);
  #10;

  //CASE: 100
  SFN=2'b00;
  A=32'b11111110110111001011101010011000;
  B=5'b10000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(100,Y,32'b10111010100110000000000000000000);
  #10;

  //CASE: 101
  SFN=2'b01;
  A=32'b11111110110111001011101010011000;
  B=5'b10000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(101,Y,32'b00000000000000001111111011011100);
  #10;

  //CASE: 102
  SFN=2'b11;
  A=32'b11111110110111001011101010011000;
  B=5'b10000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(102,Y,32'b11111111111111111111111011011100);
  #10;

  //CASE: 103
  SFN=2'b00;
  A=32'b11111110110111001011101010011000;
  B=5'b11111;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(103,Y,32'b00000000000000000000000000000000);
  #10;

  //CASE: 104
  SFN=2'b01;
  A=32'b11111110110111001011101010011000;
  B=5'b11111;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(104,Y,32'b00000000000000000000000000000001);
  #10;

  //CASE: 105
  SFN=2'b11;
  A=32'b11111110110111001011101010011000;
  B=5'b11111;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(105,Y,32'b11111111111111111111111111111111);
  #10;


  if(weAreOk) $display("TEST OK\n\nPassed");


  end

endmodule

