`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Abdelrahman Elbehery
//
// Create Date:   01:11:09 02/10/2017
// Design Name:   REGFILE
// Module Name:   F:/Self learning/FPGA/Projects/BETA_ISE/TB_REGFILE.v
// Project Name:  BETA_ISE
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: REGFILE
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module TB_REGFILE;

  reg CLK=0;
  integer weAreOk=1;

  task PRINT;
    input integer CN;
    input [31:0] RADATA;
    input [31:0] ExRADATA;
    input [31:0] RBDATA;
    input [31:0] ExRBDATA;
    if( RADATA!=ExRADATA | RBDATA!=ExRBDATA ) begin
    $display("Error in case: %d\nRADATA: %b\nExpected: %b\nRBDATA: %b\nExpected: %b\n",CN,RADATA,ExRADATA,RBDATA,ExRBDATA);
    weAreOk=0;
    end
  endtask

  reg  RA2SEL;
  reg  WASEL;
  reg  WERF;
  reg [4:0] RA;
  reg [4:0] RB;
  reg [4:0] RC;
  reg [31:0] WDATA;
  wire [31:0] RADATA;
  wire [31:0] RBDATA;

  REGFILE uut(.CLK(CLK),.RA2SEL(RA2SEL),.WASEL(WASEL),.WERF(WERF),.RA(RA),.RB(RB),.RC(RC),.WDATA(WDATA),.RADATA(RADATA),.RBDATA(RBDATA));



initial begin
  //CASE: 1
  RA2SEL=1'b0;
  WASEL=1'b0;
  WERF=1'b0;
  RA=5'b11111;
  RB=5'b11111;
  RC=5'b00000;
  WDATA=32'b00000000000000000000000000000000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(1,RADATA,32'b00000000000000000000000000000000,RBDATA,32'b00000000000000000000000000000000);
  #10;

  //CASE: 2
  RA2SEL=1'b0;
  WASEL=1'b0;
  WERF=1'b1;
  RA=5'b00000;
  RB=5'b00000;
  RC=5'b00000;
  WDATA=32'b00000000000000000000000000000000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(2,RADATA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx,RBDATA,32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
  #10;

  //CASE: 3
  RA2SEL=1'b0;
  WASEL=1'b0;
  WERF=1'b1;
  RA=5'b00000;
  RB=5'b00000;
  RC=5'b00001;
  WDATA=32'b00000000000000000000000000000001;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(3,RADATA,32'b00000000000000000000000000000000,RBDATA,32'b00000000000000000000000000000000);
  #10;

  //CASE: 4
  RA2SEL=1'b0;
  WASEL=1'b0;
  WERF=1'b1;
  RA=5'b00001;
  RB=5'b00000;
  RC=5'b00010;
  WDATA=32'b00000000000000000000000000000010;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(4,RADATA,32'b00000000000000000000000000000001,RBDATA,32'b00000000000000000000000000000000);
  #10;

  //CASE: 5
  RA2SEL=1'b0;
  WASEL=1'b0;
  WERF=1'b1;
  RA=5'b00010;
  RB=5'b00001;
  RC=5'b00011;
  WDATA=32'b00000000000000000000000000000011;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(5,RADATA,32'b00000000000000000000000000000010,RBDATA,32'b00000000000000000000000000000001);
  #10;

  //CASE: 6
  RA2SEL=1'b0;
  WASEL=1'b0;
  WERF=1'b1;
  RA=5'b00011;
  RB=5'b00010;
  RC=5'b00100;
  WDATA=32'b00000000000000000000000000000100;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(6,RADATA,32'b00000000000000000000000000000011,RBDATA,32'b00000000000000000000000000000010);
  #10;

  //CASE: 7
  RA2SEL=1'b0;
  WASEL=1'b0;
  WERF=1'b1;
  RA=5'b00100;
  RB=5'b00011;
  RC=5'b00101;
  WDATA=32'b00000000000000000000000000000101;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(7,RADATA,32'b00000000000000000000000000000100,RBDATA,32'b00000000000000000000000000000011);
  #10;

  //CASE: 8
  RA2SEL=1'b0;
  WASEL=1'b0;
  WERF=1'b1;
  RA=5'b00101;
  RB=5'b00100;
  RC=5'b00110;
  WDATA=32'b00000000000000000000000000000110;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(8,RADATA,32'b00000000000000000000000000000101,RBDATA,32'b00000000000000000000000000000100);
  #10;

  //CASE: 9
  RA2SEL=1'b0;
  WASEL=1'b0;
  WERF=1'b1;
  RA=5'b00110;
  RB=5'b00101;
  RC=5'b00111;
  WDATA=32'b00000000000000000000000000000111;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(9,RADATA,32'b00000000000000000000000000000110,RBDATA,32'b00000000000000000000000000000101);
  #10;

  //CASE: 10
  RA2SEL=1'b0;
  WASEL=1'b0;
  WERF=1'b1;
  RA=5'b00111;
  RB=5'b00110;
  RC=5'b01000;
  WDATA=32'b00000000000000000000000000001000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(10,RADATA,32'b00000000000000000000000000000111,RBDATA,32'b00000000000000000000000000000110);
  #10;

  //CASE: 11
  RA2SEL=1'b0;
  WASEL=1'b0;
  WERF=1'b1;
  RA=5'b01000;
  RB=5'b00111;
  RC=5'b01001;
  WDATA=32'b00000000000000000000000000001001;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(11,RADATA,32'b00000000000000000000000000001000,RBDATA,32'b00000000000000000000000000000111);
  #10;

  //CASE: 12
  RA2SEL=1'b0;
  WASEL=1'b0;
  WERF=1'b1;
  RA=5'b01001;
  RB=5'b01000;
  RC=5'b01010;
  WDATA=32'b00000000000000000000000000001010;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(12,RADATA,32'b00000000000000000000000000001001,RBDATA,32'b00000000000000000000000000001000);
  #10;

  //CASE: 13
  RA2SEL=1'b0;
  WASEL=1'b0;
  WERF=1'b1;
  RA=5'b01010;
  RB=5'b01001;
  RC=5'b01011;
  WDATA=32'b00000000000000000000000000001011;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(13,RADATA,32'b00000000000000000000000000001010,RBDATA,32'b00000000000000000000000000001001);
  #10;

  //CASE: 14
  RA2SEL=1'b0;
  WASEL=1'b0;
  WERF=1'b1;
  RA=5'b01011;
  RB=5'b01010;
  RC=5'b01100;
  WDATA=32'b00000000000000000000000000001100;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(14,RADATA,32'b00000000000000000000000000001011,RBDATA,32'b00000000000000000000000000001010);
  #10;

  //CASE: 15
  RA2SEL=1'b0;
  WASEL=1'b0;
  WERF=1'b1;
  RA=5'b01100;
  RB=5'b01011;
  RC=5'b01101;
  WDATA=32'b00000000000000000000000000001101;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(15,RADATA,32'b00000000000000000000000000001100,RBDATA,32'b00000000000000000000000000001011);
  #10;

  //CASE: 16
  RA2SEL=1'b0;
  WASEL=1'b0;
  WERF=1'b1;
  RA=5'b01101;
  RB=5'b01100;
  RC=5'b01110;
  WDATA=32'b00000000000000000000000000001110;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(16,RADATA,32'b00000000000000000000000000001101,RBDATA,32'b00000000000000000000000000001100);
  #10;

  //CASE: 17
  RA2SEL=1'b0;
  WASEL=1'b0;
  WERF=1'b1;
  RA=5'b01110;
  RB=5'b01101;
  RC=5'b01111;
  WDATA=32'b00000000000000000000000000001111;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(17,RADATA,32'b00000000000000000000000000001110,RBDATA,32'b00000000000000000000000000001101);
  #10;

  //CASE: 18
  RA2SEL=1'b0;
  WASEL=1'b0;
  WERF=1'b1;
  RA=5'b01111;
  RB=5'b01110;
  RC=5'b10000;
  WDATA=32'b00000000000000000000000000010000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(18,RADATA,32'b00000000000000000000000000001111,RBDATA,32'b00000000000000000000000000001110);
  #10;

  //CASE: 19
  RA2SEL=1'b0;
  WASEL=1'b0;
  WERF=1'b1;
  RA=5'b10000;
  RB=5'b01111;
  RC=5'b10001;
  WDATA=32'b00000000000000000000000000010001;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(19,RADATA,32'b00000000000000000000000000010000,RBDATA,32'b00000000000000000000000000001111);
  #10;

  //CASE: 20
  RA2SEL=1'b0;
  WASEL=1'b0;
  WERF=1'b1;
  RA=5'b10001;
  RB=5'b10000;
  RC=5'b10010;
  WDATA=32'b00000000000000000000000000010010;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(20,RADATA,32'b00000000000000000000000000010001,RBDATA,32'b00000000000000000000000000010000);
  #10;

  //CASE: 21
  RA2SEL=1'b0;
  WASEL=1'b0;
  WERF=1'b1;
  RA=5'b10010;
  RB=5'b10001;
  RC=5'b10011;
  WDATA=32'b00000000000000000000000000010011;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(21,RADATA,32'b00000000000000000000000000010010,RBDATA,32'b00000000000000000000000000010001);
  #10;

  //CASE: 22
  RA2SEL=1'b0;
  WASEL=1'b0;
  WERF=1'b1;
  RA=5'b10011;
  RB=5'b10010;
  RC=5'b10100;
  WDATA=32'b00000000000000000000000000010100;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(22,RADATA,32'b00000000000000000000000000010011,RBDATA,32'b00000000000000000000000000010010);
  #10;

  //CASE: 23
  RA2SEL=1'b0;
  WASEL=1'b0;
  WERF=1'b1;
  RA=5'b10100;
  RB=5'b10011;
  RC=5'b10101;
  WDATA=32'b00000000000000000000000000010101;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(23,RADATA,32'b00000000000000000000000000010100,RBDATA,32'b00000000000000000000000000010011);
  #10;

  //CASE: 24
  RA2SEL=1'b0;
  WASEL=1'b0;
  WERF=1'b1;
  RA=5'b10101;
  RB=5'b10100;
  RC=5'b10110;
  WDATA=32'b00000000000000000000000000010110;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(24,RADATA,32'b00000000000000000000000000010101,RBDATA,32'b00000000000000000000000000010100);
  #10;

  //CASE: 25
  RA2SEL=1'b0;
  WASEL=1'b0;
  WERF=1'b1;
  RA=5'b10110;
  RB=5'b10101;
  RC=5'b10111;
  WDATA=32'b00000000000000000000000000010111;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(25,RADATA,32'b00000000000000000000000000010110,RBDATA,32'b00000000000000000000000000010101);
  #10;

  //CASE: 26
  RA2SEL=1'b0;
  WASEL=1'b0;
  WERF=1'b1;
  RA=5'b10111;
  RB=5'b10110;
  RC=5'b11000;
  WDATA=32'b00000000000000000000000000011000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(26,RADATA,32'b00000000000000000000000000010111,RBDATA,32'b00000000000000000000000000010110);
  #10;

  //CASE: 27
  RA2SEL=1'b0;
  WASEL=1'b0;
  WERF=1'b1;
  RA=5'b11000;
  RB=5'b10111;
  RC=5'b11001;
  WDATA=32'b00000000000000000000000000011001;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(27,RADATA,32'b00000000000000000000000000011000,RBDATA,32'b00000000000000000000000000010111);
  #10;

  //CASE: 28
  RA2SEL=1'b0;
  WASEL=1'b0;
  WERF=1'b1;
  RA=5'b11001;
  RB=5'b11000;
  RC=5'b11010;
  WDATA=32'b00000000000000000000000000011010;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(28,RADATA,32'b00000000000000000000000000011001,RBDATA,32'b00000000000000000000000000011000);
  #10;

  //CASE: 29
  RA2SEL=1'b0;
  WASEL=1'b0;
  WERF=1'b1;
  RA=5'b11010;
  RB=5'b11001;
  RC=5'b11011;
  WDATA=32'b00000000000000000000000000011011;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(29,RADATA,32'b00000000000000000000000000011010,RBDATA,32'b00000000000000000000000000011001);
  #10;

  //CASE: 30
  RA2SEL=1'b0;
  WASEL=1'b0;
  WERF=1'b1;
  RA=5'b11011;
  RB=5'b11010;
  RC=5'b11100;
  WDATA=32'b00000000000000000000000000011100;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(30,RADATA,32'b00000000000000000000000000011011,RBDATA,32'b00000000000000000000000000011010);
  #10;

  //CASE: 31
  RA2SEL=1'b0;
  WASEL=1'b0;
  WERF=1'b1;
  RA=5'b11100;
  RB=5'b11011;
  RC=5'b11101;
  WDATA=32'b00000000000000000000000000011101;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(31,RADATA,32'b00000000000000000000000000011100,RBDATA,32'b00000000000000000000000000011011);
  #10;

  //CASE: 32
  RA2SEL=1'b0;
  WASEL=1'b0;
  WERF=1'b1;
  RA=5'b11101;
  RB=5'b11100;
  RC=5'b11110;
  WDATA=32'b00000000000000000000000000011110;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(32,RADATA,32'b00000000000000000000000000011101,RBDATA,32'b00000000000000000000000000011100);
  #10;

  //CASE: 33
  RA2SEL=1'b0;
  WASEL=1'b0;
  WERF=1'b1;
  RA=5'b11110;
  RB=5'b11101;
  RC=5'b11111;
  WDATA=32'b00000000000000000000000000011111;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(33,RADATA,32'b00000000000000000000000000011110,RBDATA,32'b00000000000000000000000000011101);
  #10;

  //CASE: 34
  RA2SEL=1'b0;
  WASEL=1'b0;
  WERF=1'b0;
  RA=5'b11111;
  RB=5'b11110;
  RC=5'b11111;
  WDATA=32'b00000000000000000000000000000000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(34,RADATA,32'b00000000000000000000000000000000,RBDATA,32'b00000000000000000000000000011110);
  #10;

  //CASE: 35
  RA2SEL=1'b0;
  WASEL=1'b0;
  WERF=1'b0;
  RA=5'b00000;
  RB=5'b11111;
  RC=5'b11111;
  WDATA=32'b00000000000000000000000000000000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(35,RADATA,32'b00000000000000000000000000000000,RBDATA,32'b00000000000000000000000000000000);
  #10;

  //CASE: 36
  RA2SEL=1'b1;
  WASEL=1'b0;
  WERF=1'b0;
  RA=5'b00001;
  RB=5'b00010;
  RC=5'b00011;
  WDATA=32'b00000000000000000000000000000000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(36,RADATA,32'b00000000000000000000000000000001,RBDATA,32'b00000000000000000000000000000011);
  #10;

  //CASE: 37
  RA2SEL=1'b1;
  WASEL=1'b0;
  WERF=1'b0;
  RA=5'b00001;
  RB=5'b00010;
  RC=5'b11111;
  WDATA=32'b00000000000000000000000000000000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(37,RADATA,32'b00000000000000000000000000000001,RBDATA,32'b00000000000000000000000000000000);
  #10;

  //CASE: 38
  RA2SEL=1'b1;
  WASEL=1'b0;
  WERF=1'b0;
  RA=5'b00001;
  RB=5'b11111;
  RC=5'b00100;
  WDATA=32'b00000000000000000000000000000000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(38,RADATA,32'b00000000000000000000000000000001,RBDATA,32'b00000000000000000000000000000100);
  #10;

  //CASE: 39
  RA2SEL=1'b0;
  WASEL=1'b1;
  WERF=1'b1;
  RA=5'b00001;
  RB=5'b00010;
  RC=5'b11111;
  WDATA=32'b00000000000000000011000000111001;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(39,RADATA,32'b00000000000000000000000000000001,RBDATA,32'b00000000000000000000000000000010);
  #10;

  //CASE: 40
  RA2SEL=1'b0;
  WASEL=1'b0;
  WERF=1'b0;
  RA=5'b11110;
  RB=5'b00001;
  RC=5'b00010;
  WDATA=32'b00000000000000000000000000000000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(40,RADATA,32'b00000000000000000011000000111001,RBDATA,32'b00000000000000000000000000000001);
  #10;

  //CASE: 41
  RA2SEL=1'b0;
  WASEL=1'b1;
  WERF=1'b1;
  RA=5'b00001;
  RB=5'b00010;
  RC=5'b00011;
  WDATA=32'b00000000101111000110000101001110;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(41,RADATA,32'b00000000000000000000000000000001,RBDATA,32'b00000000000000000000000000000010);
  #10;

  //CASE: 42
  RA2SEL=1'b1;
  WASEL=1'b0;
  WERF=1'b0;
  RA=5'b11110;
  RB=5'b00010;
  RC=5'b11110;
  WDATA=32'b00000000000000000000000000000000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(42,RADATA,32'b00000000101111000110000101001110,RBDATA,32'b00000000101111000110000101001110);
  #10;

  //CASE: 43
  RA2SEL=1'b0;
  WASEL=1'b0;
  WERF=1'b0;
  RA=5'b00001;
  RB=5'b00010;
  RC=5'b00011;
  WDATA=32'b00000000101111000110000101001110;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(43,RADATA,32'b00000000000000000000000000000001,RBDATA,32'b00000000000000000000000000000010);
  #10;

  //CASE: 44
  RA2SEL=1'b0;
  WASEL=1'b0;
  WERF=1'b0;
  RA=5'b00011;
  RB=5'b00011;
  RC=5'b00011;
  WDATA=32'b00000000101111000110000101001110;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(44,RADATA,32'b00000000000000000000000000000011,RBDATA,32'b00000000000000000000000000000011);
  #10;


  if(weAreOk) $display("TEST OK\n\nPassed");
  
//  RA=1;
//  #1;
//  CLK=1;#1;CLK=0;#1;
  end

endmodule