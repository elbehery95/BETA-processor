`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Abdelrahman Elbehery
//
// Create Date:   00:19:58 02/10/2017
// Design Name:   ALU
// Module Name:   F:/Self learning/FPGA/Projects/BETA_ISE/TB_ALU.v
// Project Name:  BETA_ISE
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: ALU
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module TB_ALU;

  reg CLK=0;
  integer weAreOk=1;

  task PRINT;
    input integer CN;
    input [31:0] Y;
    input [31:0] ExY;
  input Z;
  input ExZ;
  input V;
  input ExV;
  input N;
  input ExN;
    if( Y!=ExY | Z!=ExZ | V!=ExV | N!=ExN ) begin
    $display("Error in case: %d\nY: %b\nExpected: %b\nZ: %b\nExpected: %b\nV: %b\nExpected: %b\nN: %b\nExpected: %b\n",CN,Y,ExY,Z,ExZ,V,ExV,N,ExN);
    weAreOk=0;
    end
  endtask

  reg [5:0] FN;
  reg [31:0] A;
  reg [31:0] B;
  wire [31:0] Y;
  wire  Z;
  wire  V;
  wire  N;

  ALU uut(.FN(FN),.A(A),.B(B),.Y(Y),.Z(Z),.V(V),.N(N));



initial begin
  //CASE: 1
  FN=6'b100000;
  A=32'b11111111000000001111111100000000;
  B=32'b11111111111111110000000000000000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(1,Y,32'b00000000000000000000000000000000,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 2
  FN=6'b100001;
  A=32'b11111111000000001111111100000000;
  B=32'b11111111111111110000000000000000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(2,Y,32'b00000000000000000000000011111111,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 3
  FN=6'b100010;
  A=32'b11111111000000001111111100000000;
  B=32'b11111111111111110000000000000000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(3,Y,32'b00000000000000001111111100000000,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 4
  FN=6'b100011;
  A=32'b11111111000000001111111100000000;
  B=32'b11111111111111110000000000000000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(4,Y,32'b00000000000000001111111111111111,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 5
  FN=6'b100100;
  A=32'b11111111000000001111111100000000;
  B=32'b11111111111111110000000000000000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(5,Y,32'b00000000111111110000000000000000,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 6
  FN=6'b100101;
  A=32'b11111111000000001111111100000000;
  B=32'b11111111111111110000000000000000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(6,Y,32'b00000000111111110000000011111111,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 7
  FN=6'b100110;
  A=32'b11111111000000001111111100000000;
  B=32'b11111111111111110000000000000000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(7,Y,32'b00000000111111111111111100000000,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 8
  FN=6'b100111;
  A=32'b11111111000000001111111100000000;
  B=32'b11111111111111110000000000000000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(8,Y,32'b00000000111111111111111111111111,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 9
  FN=6'b101000;
  A=32'b11111111000000001111111100000000;
  B=32'b11111111111111110000000000000000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(9,Y,32'b11111111000000000000000000000000,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 10
  FN=6'b101001;
  A=32'b11111111000000001111111100000000;
  B=32'b11111111111111110000000000000000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(10,Y,32'b11111111000000000000000011111111,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 11
  FN=6'b101010;
  A=32'b11111111000000001111111100000000;
  B=32'b11111111111111110000000000000000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(11,Y,32'b11111111000000001111111100000000,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 12
  FN=6'b101011;
  A=32'b11111111000000001111111100000000;
  B=32'b11111111111111110000000000000000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(12,Y,32'b11111111000000001111111111111111,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 13
  FN=6'b101100;
  A=32'b11111111000000001111111100000000;
  B=32'b11111111111111110000000000000000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(13,Y,32'b11111111111111110000000000000000,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 14
  FN=6'b101101;
  A=32'b11111111000000001111111100000000;
  B=32'b11111111111111110000000000000000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(14,Y,32'b11111111111111110000000011111111,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 15
  FN=6'b101110;
  A=32'b11111111000000001111111100000000;
  B=32'b11111111111111110000000000000000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(15,Y,32'b11111111111111111111111100000000,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 16
  FN=6'b101111;
  A=32'b11111111000000001111111100000000;
  B=32'b11111111111111110000000000000000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(16,Y,32'b11111111111111111111111111111111,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 17
  FN=6'b110000;
  A=32'b00000000000000000000000000000000;
  B=32'b00000000000000000000000000000000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(17,Y,32'b00000000000000000000000000000000,Z,1'b1,V,1'b0,N,1'b0);
  #10;

  //CASE: 18
  FN=6'b110001;
  A=32'b00000000000000000000000000000000;
  B=32'b00000000000000000000000000000000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(18,Y,32'b00000000000000000000000000000000,Z,1'b1,V,1'b0,N,1'b0);
  #10;

  //CASE: 19
  FN=6'b110011;
  A=32'b00000000000000000000000000000000;
  B=32'b00000000000000000000000000000000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(19,Y,32'b00000000000000000000000000000000,Z,1'b1,V,1'b0,N,1'b0);
  #10;

  //CASE: 20
  FN=6'b110000;
  A=32'b00000000000000000000000000000000;
  B=32'b00000000000000000000000000000001;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(20,Y,32'b00000000000000000000000000000000,Z,1'b0,V,1'b0,N,1'b0);
  #10;

  //CASE: 21
  FN=6'b110001;
  A=32'b00000000000000000000000000000000;
  B=32'b00000000000000000000000000000001;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(21,Y,32'b00000000000000000000000000000000,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 22
  FN=6'b110011;
  A=32'b00000000000000000000000000000000;
  B=32'b00000000000000000000000000000001;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(22,Y,32'b00000000000000000000000000000000,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 23
  FN=6'b110000;
  A=32'b00000000000000000000000000000000;
  B=32'b00000000000000000000000000000010;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(23,Y,32'b00000000000000000000000000000000,Z,1'b0,V,1'b0,N,1'b0);
  #10;

  //CASE: 24
  FN=6'b110001;
  A=32'b00000000000000000000000000000000;
  B=32'b00000000000000000000000000000010;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(24,Y,32'b00000000000000000000000000000000,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 25
  FN=6'b110011;
  A=32'b00000000000000000000000000000000;
  B=32'b00000000000000000000000000000010;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(25,Y,32'b00000000000000000000000000000000,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 26
  FN=6'b110000;
  A=32'b00000000000000000000000000000000;
  B=32'b00000000000000000000000000000100;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(26,Y,32'b00000000000000000000000000000000,Z,1'b0,V,1'b0,N,1'b0);
  #10;

  //CASE: 27
  FN=6'b110001;
  A=32'b00000000000000000000000000000000;
  B=32'b00000000000000000000000000000100;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(27,Y,32'b00000000000000000000000000000000,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 28
  FN=6'b110011;
  A=32'b00000000000000000000000000000000;
  B=32'b00000000000000000000000000000100;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(28,Y,32'b00000000000000000000000000000000,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 29
  FN=6'b110000;
  A=32'b00000000000000000000000000000000;
  B=32'b00000000000000000000000000001000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(29,Y,32'b00000000000000000000000000000000,Z,1'b0,V,1'b0,N,1'b0);
  #10;

  //CASE: 30
  FN=6'b110001;
  A=32'b00000000000000000000000000000000;
  B=32'b00000000000000000000000000001000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(30,Y,32'b00000000000000000000000000000000,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 31
  FN=6'b110011;
  A=32'b00000000000000000000000000000000;
  B=32'b00000000000000000000000000001000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(31,Y,32'b00000000000000000000000000000000,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 32
  FN=6'b110000;
  A=32'b00000000000000000000000000000000;
  B=32'b00000000000000000000000000010000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(32,Y,32'b00000000000000000000000000000000,Z,1'b0,V,1'b0,N,1'b0);
  #10;

  //CASE: 33
  FN=6'b110001;
  A=32'b00000000000000000000000000000000;
  B=32'b00000000000000000000000000010000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(33,Y,32'b00000000000000000000000000000000,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 34
  FN=6'b110011;
  A=32'b00000000000000000000000000000000;
  B=32'b00000000000000000000000000010000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(34,Y,32'b00000000000000000000000000000000,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 35
  FN=6'b110000;
  A=32'b00000000000000000000000000000000;
  B=32'b00000000000000000000000000011111;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(35,Y,32'b00000000000000000000000000000000,Z,1'b0,V,1'b0,N,1'b0);
  #10;

  //CASE: 36
  FN=6'b110001;
  A=32'b00000000000000000000000000000000;
  B=32'b00000000000000000000000000011111;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(36,Y,32'b00000000000000000000000000000000,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 37
  FN=6'b110011;
  A=32'b00000000000000000000000000000000;
  B=32'b00000000000000000000000000011111;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(37,Y,32'b00000000000000000000000000000000,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 38
  FN=6'b110000;
  A=32'b00000000000000000000000000000001;
  B=32'b00000000000000000000000000000000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(38,Y,32'b00000000000000000000000000000001,Z,1'b0,V,1'b0,N,1'b0);
  #10;

  //CASE: 39
  FN=6'b110001;
  A=32'b00000000000000000000000000000001;
  B=32'b00000000000000000000000000000000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(39,Y,32'b00000000000000000000000000000001,Z,1'b0,V,1'b0,N,1'b0);
  #10;

  //CASE: 40
  FN=6'b110011;
  A=32'b00000000000000000000000000000001;
  B=32'b00000000000000000000000000000000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(40,Y,32'b00000000000000000000000000000001,Z,1'b0,V,1'b0,N,1'b0);
  #10;

  //CASE: 41
  FN=6'b110000;
  A=32'b00000000000000000000000000000001;
  B=32'b00000000000000000000000000000001;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(41,Y,32'b00000000000000000000000000000010,Z,1'b0,V,1'b0,N,1'b0);
  #10;

  //CASE: 42
  FN=6'b110001;
  A=32'b00000000000000000000000000000001;
  B=32'b00000000000000000000000000000001;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(42,Y,32'b00000000000000000000000000000000,Z,1'b1,V,1'b0,N,1'b0);
  #10;

  //CASE: 43
  FN=6'b110011;
  A=32'b00000000000000000000000000000001;
  B=32'b00000000000000000000000000000001;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(43,Y,32'b00000000000000000000000000000000,Z,1'b1,V,1'b0,N,1'b0);
  #10;

  //CASE: 44
  FN=6'b110000;
  A=32'b00000000000000000000000000000001;
  B=32'b00000000000000000000000000000010;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(44,Y,32'b00000000000000000000000000000100,Z,1'b0,V,1'b0,N,1'b0);
  #10;

  //CASE: 45
  FN=6'b110001;
  A=32'b00000000000000000000000000000001;
  B=32'b00000000000000000000000000000010;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(45,Y,32'b00000000000000000000000000000000,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 46
  FN=6'b110011;
  A=32'b00000000000000000000000000000001;
  B=32'b00000000000000000000000000000010;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(46,Y,32'b00000000000000000000000000000000,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 47
  FN=6'b110000;
  A=32'b00000000000000000000000000000001;
  B=32'b00000000000000000000000000000100;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(47,Y,32'b00000000000000000000000000010000,Z,1'b0,V,1'b0,N,1'b0);
  #10;

  //CASE: 48
  FN=6'b110001;
  A=32'b00000000000000000000000000000001;
  B=32'b00000000000000000000000000000100;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(48,Y,32'b00000000000000000000000000000000,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 49
  FN=6'b110011;
  A=32'b00000000000000000000000000000001;
  B=32'b00000000000000000000000000000100;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(49,Y,32'b00000000000000000000000000000000,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 50
  FN=6'b110000;
  A=32'b00000000000000000000000000000001;
  B=32'b00000000000000000000000000001000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(50,Y,32'b00000000000000000000000100000000,Z,1'b0,V,1'b0,N,1'b0);
  #10;

  //CASE: 51
  FN=6'b110001;
  A=32'b00000000000000000000000000000001;
  B=32'b00000000000000000000000000001000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(51,Y,32'b00000000000000000000000000000000,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 52
  FN=6'b110011;
  A=32'b00000000000000000000000000000001;
  B=32'b00000000000000000000000000001000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(52,Y,32'b00000000000000000000000000000000,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 53
  FN=6'b110000;
  A=32'b00000000000000000000000000000001;
  B=32'b00000000000000000000000000010000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(53,Y,32'b00000000000000010000000000000000,Z,1'b0,V,1'b0,N,1'b0);
  #10;

  //CASE: 54
  FN=6'b110001;
  A=32'b00000000000000000000000000000001;
  B=32'b00000000000000000000000000010000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(54,Y,32'b00000000000000000000000000000000,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 55
  FN=6'b110011;
  A=32'b00000000000000000000000000000001;
  B=32'b00000000000000000000000000010000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(55,Y,32'b00000000000000000000000000000000,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 56
  FN=6'b110000;
  A=32'b00000000000000000000000000000001;
  B=32'b00000000000000000000000000011111;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(56,Y,32'b10000000000000000000000000000000,Z,1'b0,V,1'b0,N,1'b0);
  #10;

  //CASE: 57
  FN=6'b110001;
  A=32'b00000000000000000000000000000001;
  B=32'b00000000000000000000000000011111;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(57,Y,32'b00000000000000000000000000000000,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 58
  FN=6'b110011;
  A=32'b00000000000000000000000000000001;
  B=32'b00000000000000000000000000011111;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(58,Y,32'b00000000000000000000000000000000,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 59
  FN=6'b110000;
  A=32'b11111111111111111111111111111111;
  B=32'b00000000000000000000000000000000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(59,Y,32'b11111111111111111111111111111111,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 60
  FN=6'b110001;
  A=32'b11111111111111111111111111111111;
  B=32'b00000000000000000000000000000000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(60,Y,32'b11111111111111111111111111111111,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 61
  FN=6'b110011;
  A=32'b11111111111111111111111111111111;
  B=32'b00000000000000000000000000000000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(61,Y,32'b11111111111111111111111111111111,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 62
  FN=6'b110000;
  A=32'b11111111111111111111111111111111;
  B=32'b00000000000000000000000000000001;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(62,Y,32'b11111111111111111111111111111110,Z,1'b1,V,1'b0,N,1'b0);
  #10;

  //CASE: 63
  FN=6'b110001;
  A=32'b11111111111111111111111111111111;
  B=32'b00000000000000000000000000000001;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(63,Y,32'b01111111111111111111111111111111,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 64
  FN=6'b110011;
  A=32'b11111111111111111111111111111111;
  B=32'b00000000000000000000000000000001;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(64,Y,32'b11111111111111111111111111111111,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 65
  FN=6'b110000;
  A=32'b11111111111111111111111111111111;
  B=32'b00000000000000000000000000000010;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(65,Y,32'b11111111111111111111111111111100,Z,1'b0,V,1'b0,N,1'b0);
  #10;

  //CASE: 66
  FN=6'b110001;
  A=32'b11111111111111111111111111111111;
  B=32'b00000000000000000000000000000010;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(66,Y,32'b00111111111111111111111111111111,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 67
  FN=6'b110011;
  A=32'b11111111111111111111111111111111;
  B=32'b00000000000000000000000000000010;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(67,Y,32'b11111111111111111111111111111111,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 68
  FN=6'b110000;
  A=32'b11111111111111111111111111111111;
  B=32'b00000000000000000000000000000100;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(68,Y,32'b11111111111111111111111111110000,Z,1'b0,V,1'b0,N,1'b0);
  #10;

  //CASE: 69
  FN=6'b110001;
  A=32'b11111111111111111111111111111111;
  B=32'b00000000000000000000000000000100;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(69,Y,32'b00001111111111111111111111111111,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 70
  FN=6'b110011;
  A=32'b11111111111111111111111111111111;
  B=32'b00000000000000000000000000000100;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(70,Y,32'b11111111111111111111111111111111,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 71
  FN=6'b110000;
  A=32'b11111111111111111111111111111111;
  B=32'b00000000000000000000000000001000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(71,Y,32'b11111111111111111111111100000000,Z,1'b0,V,1'b0,N,1'b0);
  #10;

  //CASE: 72
  FN=6'b110001;
  A=32'b11111111111111111111111111111111;
  B=32'b00000000000000000000000000001000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(72,Y,32'b00000000111111111111111111111111,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 73
  FN=6'b110011;
  A=32'b11111111111111111111111111111111;
  B=32'b00000000000000000000000000001000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(73,Y,32'b11111111111111111111111111111111,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 74
  FN=6'b110000;
  A=32'b11111111111111111111111111111111;
  B=32'b00000000000000000000000000010000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(74,Y,32'b11111111111111110000000000000000,Z,1'b0,V,1'b0,N,1'b0);
  #10;

  //CASE: 75
  FN=6'b110001;
  A=32'b11111111111111111111111111111111;
  B=32'b00000000000000000000000000010000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(75,Y,32'b00000000000000001111111111111111,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 76
  FN=6'b110011;
  A=32'b11111111111111111111111111111111;
  B=32'b00000000000000000000000000010000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(76,Y,32'b11111111111111111111111111111111,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 77
  FN=6'b110000;
  A=32'b11111111111111111111111111111111;
  B=32'b00000000000000000000000000011111;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(77,Y,32'b10000000000000000000000000000000,Z,1'b0,V,1'b0,N,1'b0);
  #10;

  //CASE: 78
  FN=6'b110001;
  A=32'b11111111111111111111111111111111;
  B=32'b00000000000000000000000000011111;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(78,Y,32'b00000000000000000000000000000001,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 79
  FN=6'b110011;
  A=32'b11111111111111111111111111111111;
  B=32'b00000000000000000000000000011111;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(79,Y,32'b11111111111111111111111111111111,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 80
  FN=6'b110000;
  A=32'b00010010001101000101011001111000;
  B=32'b00000000000000000000000000000000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(80,Y,32'b00010010001101000101011001111000,Z,1'b0,V,1'b0,N,1'b0);
  #10;

  //CASE: 81
  FN=6'b110001;
  A=32'b00010010001101000101011001111000;
  B=32'b00000000000000000000000000000000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(81,Y,32'b00010010001101000101011001111000,Z,1'b0,V,1'b0,N,1'b0);
  #10;

  //CASE: 82
  FN=6'b110011;
  A=32'b00010010001101000101011001111000;
  B=32'b00000000000000000000000000000000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(82,Y,32'b00010010001101000101011001111000,Z,1'b0,V,1'b0,N,1'b0);
  #10;

  //CASE: 83
  FN=6'b110000;
  A=32'b00010010001101000101011001111000;
  B=32'b00000000000000000000000000000001;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(83,Y,32'b00100100011010001010110011110000,Z,1'b0,V,1'b0,N,1'b0);
  #10;

  //CASE: 84
  FN=6'b110001;
  A=32'b00010010001101000101011001111000;
  B=32'b00000000000000000000000000000001;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(84,Y,32'b00001001000110100010101100111100,Z,1'b0,V,1'b0,N,1'b0);
  #10;

  //CASE: 85
  FN=6'b110011;
  A=32'b00010010001101000101011001111000;
  B=32'b00000000000000000000000000000001;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(85,Y,32'b00001001000110100010101100111100,Z,1'b0,V,1'b0,N,1'b0);
  #10;

  //CASE: 86
  FN=6'b110000;
  A=32'b00010010001101000101011001111000;
  B=32'b00000000000000000000000000000010;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(86,Y,32'b01001000110100010101100111100000,Z,1'b0,V,1'b0,N,1'b0);
  #10;

  //CASE: 87
  FN=6'b110001;
  A=32'b00010010001101000101011001111000;
  B=32'b00000000000000000000000000000010;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(87,Y,32'b00000100100011010001010110011110,Z,1'b0,V,1'b0,N,1'b0);
  #10;

  //CASE: 88
  FN=6'b110011;
  A=32'b00010010001101000101011001111000;
  B=32'b00000000000000000000000000000010;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(88,Y,32'b00000100100011010001010110011110,Z,1'b0,V,1'b0,N,1'b0);
  #10;

  //CASE: 89
  FN=6'b110000;
  A=32'b00010010001101000101011001111000;
  B=32'b00000000000000000000000000000100;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(89,Y,32'b00100011010001010110011110000000,Z,1'b0,V,1'b0,N,1'b0);
  #10;

  //CASE: 90
  FN=6'b110001;
  A=32'b00010010001101000101011001111000;
  B=32'b00000000000000000000000000000100;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(90,Y,32'b00000001001000110100010101100111,Z,1'b0,V,1'b0,N,1'b0);
  #10;

  //CASE: 91
  FN=6'b110011;
  A=32'b00010010001101000101011001111000;
  B=32'b00000000000000000000000000000100;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(91,Y,32'b00000001001000110100010101100111,Z,1'b0,V,1'b0,N,1'b0);
  #10;

  //CASE: 92
  FN=6'b110000;
  A=32'b00010010001101000101011001111000;
  B=32'b00000000000000000000000000001000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(92,Y,32'b00110100010101100111100000000000,Z,1'b0,V,1'b0,N,1'b0);
  #10;

  //CASE: 93
  FN=6'b110001;
  A=32'b00010010001101000101011001111000;
  B=32'b00000000000000000000000000001000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(93,Y,32'b00000000000100100011010001010110,Z,1'b0,V,1'b0,N,1'b0);
  #10;

  //CASE: 94
  FN=6'b110011;
  A=32'b00010010001101000101011001111000;
  B=32'b00000000000000000000000000001000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(94,Y,32'b00000000000100100011010001010110,Z,1'b0,V,1'b0,N,1'b0);
  #10;

  //CASE: 95
  FN=6'b110000;
  A=32'b00010010001101000101011001111000;
  B=32'b00000000000000000000000000010000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(95,Y,32'b01010110011110000000000000000000,Z,1'b0,V,1'b0,N,1'b0);
  #10;

  //CASE: 96
  FN=6'b110001;
  A=32'b00010010001101000101011001111000;
  B=32'b00000000000000000000000000010000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(96,Y,32'b00000000000000000001001000110100,Z,1'b0,V,1'b0,N,1'b0);
  #10;

  //CASE: 97
  FN=6'b110011;
  A=32'b00010010001101000101011001111000;
  B=32'b00000000000000000000000000010000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(97,Y,32'b00000000000000000001001000110100,Z,1'b0,V,1'b0,N,1'b0);
  #10;

  //CASE: 98
  FN=6'b110000;
  A=32'b00010010001101000101011001111000;
  B=32'b00000000000000000000000000011111;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(98,Y,32'b00000000000000000000000000000000,Z,1'b0,V,1'b0,N,1'b0);
  #10;

  //CASE: 99
  FN=6'b110001;
  A=32'b00010010001101000101011001111000;
  B=32'b00000000000000000000000000011111;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(99,Y,32'b00000000000000000000000000000000,Z,1'b0,V,1'b0,N,1'b0);
  #10;

  //CASE: 100
  FN=6'b110011;
  A=32'b00010010001101000101011001111000;
  B=32'b00000000000000000000000000011111;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(100,Y,32'b00000000000000000000000000000000,Z,1'b0,V,1'b0,N,1'b0);
  #10;

  //CASE: 101
  FN=6'b110000;
  A=32'b11111110110111001010101110011000;
  B=32'b00000000000000000000000000000000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(101,Y,32'b11111110110111001010101110011000,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 102
  FN=6'b110001;
  A=32'b11111110110111001010101110011000;
  B=32'b00000000000000000000000000000000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(102,Y,32'b11111110110111001010101110011000,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 103
  FN=6'b110011;
  A=32'b11111110110111001010101110011000;
  B=32'b00000000000000000000000000000000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(103,Y,32'b11111110110111001010101110011000,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 104
  FN=6'b110000;
  A=32'b11111110110111001010101110011000;
  B=32'b00000000000000000000000000000001;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(104,Y,32'b11111101101110010101011100110000,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 105
  FN=6'b110001;
  A=32'b11111110110111001010101110011000;
  B=32'b00000000000000000000000000000001;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(105,Y,32'b01111111011011100101010111001100,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 106
  FN=6'b110011;
  A=32'b11111110110111001010101110011000;
  B=32'b00000000000000000000000000000001;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(106,Y,32'b11111111011011100101010111001100,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 107
  FN=6'b110000;
  A=32'b11111110110111001010101110011000;
  B=32'b00000000000000000000000000000010;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(107,Y,32'b11111011011100101010111001100000,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 108
  FN=6'b110001;
  A=32'b11111110110111001010101110011000;
  B=32'b00000000000000000000000000000010;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(108,Y,32'b00111111101101110010101011100110,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 109
  FN=6'b110011;
  A=32'b11111110110111001010101110011000;
  B=32'b00000000000000000000000000000010;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(109,Y,32'b11111111101101110010101011100110,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 110
  FN=6'b110000;
  A=32'b11111110110111001010101110011000;
  B=32'b00000000000000000000000000000100;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(110,Y,32'b11101101110010101011100110000000,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 111
  FN=6'b110001;
  A=32'b11111110110111001010101110011000;
  B=32'b00000000000000000000000000000100;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(111,Y,32'b00001111111011011100101010111001,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 112
  FN=6'b110011;
  A=32'b11111110110111001010101110011000;
  B=32'b00000000000000000000000000000100;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(112,Y,32'b11111111111011011100101010111001,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 113
  FN=6'b110000;
  A=32'b11111110110111001010101110011000;
  B=32'b00000000000000000000000000001000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(113,Y,32'b11011100101010111001100000000000,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 114
  FN=6'b110001;
  A=32'b11111110110111001010101110011000;
  B=32'b00000000000000000000000000001000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(114,Y,32'b00000000111111101101110010101011,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 115
  FN=6'b110011;
  A=32'b11111110110111001010101110011000;
  B=32'b00000000000000000000000000001000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(115,Y,32'b11111111111111101101110010101011,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 116
  FN=6'b110000;
  A=32'b11111110110111001010101110011000;
  B=32'b00000000000000000000000000010000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(116,Y,32'b10101011100110000000000000000000,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 117
  FN=6'b110001;
  A=32'b11111110110111001010101110011000;
  B=32'b00000000000000000000000000010000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(117,Y,32'b00000000000000001111111011011100,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 118
  FN=6'b110011;
  A=32'b11111110110111001010101110011000;
  B=32'b00000000000000000000000000010000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(118,Y,32'b11111111111111111111111011011100,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 119
  FN=6'b110000;
  A=32'b11111110110111001010101110011000;
  B=32'b00000000000000000000000000011111;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(119,Y,32'b00000000000000000000000000000000,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 120
  FN=6'b110001;
  A=32'b11111110110111001010101110011000;
  B=32'b00000000000000000000000000011111;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(120,Y,32'b00000000000000000000000000000001,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 121
  FN=6'b110011;
  A=32'b11111110110111001010101110011000;
  B=32'b00000000000000000000000000011111;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(121,Y,32'b11111111111111111111111111111111,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 122
  FN=6'b010000;
  A=32'b00000000000000000000000000000000;
  B=32'b00000000000000000000000000000000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(122,Y,32'b00000000000000000000000000000000,Z,1'b1,V,1'b0,N,1'b0);
  #10;

  //CASE: 123
  FN=6'b010000;
  A=32'b00000000000000000000000000000000;
  B=32'b00000000000000000000000000000001;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(123,Y,32'b00000000000000000000000000000001,Z,1'b0,V,1'b0,N,1'b0);
  #10;

  //CASE: 124
  FN=6'b010000;
  A=32'b00000000000000000000000000000000;
  B=32'b11111111111111111111111111111111;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(124,Y,32'b11111111111111111111111111111111,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 125
  FN=6'b010000;
  A=32'b00000000000000000000000000000000;
  B=32'b10101010101010101010101010101010;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(125,Y,32'b10101010101010101010101010101010,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 126
  FN=6'b010000;
  A=32'b00000000000000000000000000000000;
  B=32'b01010101010101010101010101010101;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(126,Y,32'b01010101010101010101010101010101,Z,1'b0,V,1'b0,N,1'b0);
  #10;

  //CASE: 127
  FN=6'b010000;
  A=32'b00000000000000000000000000000001;
  B=32'b00000000000000000000000000000000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(127,Y,32'b00000000000000000000000000000001,Z,1'b0,V,1'b0,N,1'b0);
  #10;

  //CASE: 128
  FN=6'b010000;
  A=32'b00000000000000000000000000000001;
  B=32'b00000000000000000000000000000001;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(128,Y,32'b00000000000000000000000000000010,Z,1'b0,V,1'b0,N,1'b0);
  #10;

  //CASE: 129
  FN=6'b010000;
  A=32'b00000000000000000000000000000001;
  B=32'b11111111111111111111111111111111;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(129,Y,32'b00000000000000000000000000000000,Z,1'b1,V,1'b0,N,1'b0);
  #10;

  //CASE: 130
  FN=6'b010000;
  A=32'b00000000000000000000000000000001;
  B=32'b10101010101010101010101010101010;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(130,Y,32'b10101010101010101010101010101011,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 131
  FN=6'b010000;
  A=32'b00000000000000000000000000000001;
  B=32'b01010101010101010101010101010101;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(131,Y,32'b01010101010101010101010101010110,Z,1'b0,V,1'b0,N,1'b0);
  #10;

  //CASE: 132
  FN=6'b010000;
  A=32'b11111111111111111111111111111111;
  B=32'b00000000000000000000000000000000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(132,Y,32'b11111111111111111111111111111111,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 133
  FN=6'b010000;
  A=32'b11111111111111111111111111111111;
  B=32'b00000000000000000000000000000001;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(133,Y,32'b00000000000000000000000000000000,Z,1'b1,V,1'b0,N,1'b0);
  #10;

  //CASE: 134
  FN=6'b010000;
  A=32'b11111111111111111111111111111111;
  B=32'b11111111111111111111111111111111;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(134,Y,32'b11111111111111111111111111111110,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 135
  FN=6'b010000;
  A=32'b11111111111111111111111111111111;
  B=32'b10101010101010101010101010101010;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(135,Y,32'b10101010101010101010101010101001,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 136
  FN=6'b010000;
  A=32'b11111111111111111111111111111111;
  B=32'b01010101010101010101010101010101;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(136,Y,32'b01010101010101010101010101010100,Z,1'b0,V,1'b0,N,1'b0);
  #10;

  //CASE: 137
  FN=6'b010000;
  A=32'b10101010101010101010101010101010;
  B=32'b00000000000000000000000000000000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(137,Y,32'b10101010101010101010101010101010,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 138
  FN=6'b010000;
  A=32'b10101010101010101010101010101010;
  B=32'b00000000000000000000000000000001;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(138,Y,32'b10101010101010101010101010101011,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 139
  FN=6'b010000;
  A=32'b10101010101010101010101010101010;
  B=32'b11111111111111111111111111111111;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(139,Y,32'b10101010101010101010101010101001,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 140
  FN=6'b010000;
  A=32'b10101010101010101010101010101010;
  B=32'b10101010101010101010101010101010;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(140,Y,32'b01010101010101010101010101010100,Z,1'b0,V,1'b1,N,1'b0);
  #10;

  //CASE: 141
  FN=6'b010000;
  A=32'b10101010101010101010101010101010;
  B=32'b01010101010101010101010101010101;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(141,Y,32'b11111111111111111111111111111111,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 142
  FN=6'b010000;
  A=32'b01010101010101010101010101010101;
  B=32'b00000000000000000000000000000000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(142,Y,32'b01010101010101010101010101010101,Z,1'b0,V,1'b0,N,1'b0);
  #10;

  //CASE: 143
  FN=6'b010000;
  A=32'b01010101010101010101010101010101;
  B=32'b00000000000000000000000000000001;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(143,Y,32'b01010101010101010101010101010110,Z,1'b0,V,1'b0,N,1'b0);
  #10;

  //CASE: 144
  FN=6'b010000;
  A=32'b01010101010101010101010101010101;
  B=32'b11111111111111111111111111111111;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(144,Y,32'b01010101010101010101010101010100,Z,1'b0,V,1'b0,N,1'b0);
  #10;

  //CASE: 145
  FN=6'b010000;
  A=32'b01010101010101010101010101010101;
  B=32'b10101010101010101010101010101010;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(145,Y,32'b11111111111111111111111111111111,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 146
  FN=6'b010000;
  A=32'b01010101010101010101010101010101;
  B=32'b01010101010101010101010101010101;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(146,Y,32'b10101010101010101010101010101010,Z,1'b0,V,1'b1,N,1'b1);
  #10;

  //CASE: 147
  FN=6'b010001;
  A=32'b00000000000000000000000000000000;
  B=32'b00000000000000000000000000000000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(147,Y,32'b00000000000000000000000000000000,Z,1'b1,V,1'b0,N,1'b0);
  #10;

  //CASE: 148
  FN=6'b010001;
  A=32'b00000000000000000000000000000000;
  B=32'b00000000000000000000000000000001;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(148,Y,32'b11111111111111111111111111111111,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 149
  FN=6'b010001;
  A=32'b00000000000000000000000000000000;
  B=32'b11111111111111111111111111111111;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(149,Y,32'b00000000000000000000000000000001,Z,1'b0,V,1'b0,N,1'b0);
  #10;

  //CASE: 150
  FN=6'b010001;
  A=32'b00000000000000000000000000000000;
  B=32'b10101010101010101010101010101010;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(150,Y,32'b01010101010101010101010101010110,Z,1'b0,V,1'b0,N,1'b0);
  #10;

  //CASE: 151
  FN=6'b010001;
  A=32'b00000000000000000000000000000000;
  B=32'b01010101010101010101010101010101;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(151,Y,32'b10101010101010101010101010101011,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 152
  FN=6'b010001;
  A=32'b00000000000000000000000000000001;
  B=32'b00000000000000000000000000000000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(152,Y,32'b00000000000000000000000000000001,Z,1'b0,V,1'b0,N,1'b0);
  #10;

  //CASE: 153
  FN=6'b010001;
  A=32'b00000000000000000000000000000001;
  B=32'b00000000000000000000000000000001;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(153,Y,32'b00000000000000000000000000000000,Z,1'b1,V,1'b0,N,1'b0);
  #10;

  //CASE: 154
  FN=6'b010001;
  A=32'b00000000000000000000000000000001;
  B=32'b11111111111111111111111111111111;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(154,Y,32'b00000000000000000000000000000010,Z,1'b0,V,1'b0,N,1'b0);
  #10;

  //CASE: 155
  FN=6'b010001;
  A=32'b00000000000000000000000000000001;
  B=32'b10101010101010101010101010101010;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(155,Y,32'b01010101010101010101010101010111,Z,1'b0,V,1'b0,N,1'b0);
  #10;

  //CASE: 156
  FN=6'b010001;
  A=32'b00000000000000000000000000000001;
  B=32'b01010101010101010101010101010101;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(156,Y,32'b10101010101010101010101010101100,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 157
  FN=6'b010001;
  A=32'b11111111111111111111111111111111;
  B=32'b00000000000000000000000000000000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(157,Y,32'b11111111111111111111111111111111,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 158
  FN=6'b010001;
  A=32'b11111111111111111111111111111111;
  B=32'b00000000000000000000000000000001;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(158,Y,32'b11111111111111111111111111111110,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 159
  FN=6'b010001;
  A=32'b11111111111111111111111111111111;
  B=32'b11111111111111111111111111111111;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(159,Y,32'b00000000000000000000000000000000,Z,1'b1,V,1'b0,N,1'b0);
  #10;

  //CASE: 160
  FN=6'b010001;
  A=32'b11111111111111111111111111111111;
  B=32'b10101010101010101010101010101010;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(160,Y,32'b01010101010101010101010101010101,Z,1'b0,V,1'b0,N,1'b0);
  #10;

  //CASE: 161
  FN=6'b010001;
  A=32'b11111111111111111111111111111111;
  B=32'b01010101010101010101010101010101;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(161,Y,32'b10101010101010101010101010101010,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 162
  FN=6'b010001;
  A=32'b10101010101010101010101010101010;
  B=32'b00000000000000000000000000000000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(162,Y,32'b10101010101010101010101010101010,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 163
  FN=6'b010001;
  A=32'b10101010101010101010101010101010;
  B=32'b00000000000000000000000000000001;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(163,Y,32'b10101010101010101010101010101001,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 164
  FN=6'b010001;
  A=32'b10101010101010101010101010101010;
  B=32'b11111111111111111111111111111111;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(164,Y,32'b10101010101010101010101010101011,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 165
  FN=6'b010001;
  A=32'b10101010101010101010101010101010;
  B=32'b10101010101010101010101010101010;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(165,Y,32'b00000000000000000000000000000000,Z,1'b1,V,1'b0,N,1'b0);
  #10;

  //CASE: 166
  FN=6'b010001;
  A=32'b10101010101010101010101010101010;
  B=32'b01010101010101010101010101010101;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(166,Y,32'b01010101010101010101010101010101,Z,1'b0,V,1'b1,N,1'b0);
  #10;

  //CASE: 167
  FN=6'b010001;
  A=32'b01010101010101010101010101010101;
  B=32'b00000000000000000000000000000000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(167,Y,32'b01010101010101010101010101010101,Z,1'b0,V,1'b0,N,1'b0);
  #10;

  //CASE: 168
  FN=6'b010001;
  A=32'b01010101010101010101010101010101;
  B=32'b00000000000000000000000000000001;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(168,Y,32'b01010101010101010101010101010100,Z,1'b0,V,1'b0,N,1'b0);
  #10;

  //CASE: 169
  FN=6'b010001;
  A=32'b01010101010101010101010101010101;
  B=32'b11111111111111111111111111111111;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(169,Y,32'b01010101010101010101010101010110,Z,1'b0,V,1'b0,N,1'b0);
  #10;

  //CASE: 170
  FN=6'b010001;
  A=32'b01010101010101010101010101010101;
  B=32'b10101010101010101010101010101010;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(170,Y,32'b10101010101010101010101010101011,Z,1'b0,V,1'b1,N,1'b1);
  #10;

  //CASE: 171
  FN=6'b010001;
  A=32'b01010101010101010101010101010101;
  B=32'b01010101010101010101010101010101;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(171,Y,32'b00000000000000000000000000000000,Z,1'b1,V,1'b0,N,1'b0);
  #10;

  //CASE: 172
  FN=6'b000011;
  A=32'b00000000000000000000000000000101;
  B=32'b11011110101011011011111011101111;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(172,Y,32'b00000000000000000000000000000000,Z,1'b0,V,1'b0,N,1'b0);
  #10;

  //CASE: 173
  FN=6'b000101;
  A=32'b00000000000000000000000000000101;
  B=32'b11011110101011011011111011101111;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(173,Y,32'b00000000000000000000000000000000,Z,1'b0,V,1'b0,N,1'b0);
  #10;

  //CASE: 174
  FN=6'b000111;
  A=32'b00000000000000000000000000000101;
  B=32'b11011110101011011011111011101111;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(174,Y,32'b00000000000000000000000000000000,Z,1'b0,V,1'b0,N,1'b0);
  #10;

  //CASE: 175
  FN=6'b000011;
  A=32'b00010010001101000101011001111000;
  B=32'b00010010001101000101011001111000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(175,Y,32'b00000000000000000000000000000001,Z,1'b1,V,1'b0,N,1'b0);
  #10;

  //CASE: 176
  FN=6'b000101;
  A=32'b00010010001101000101011001111000;
  B=32'b00010010001101000101011001111000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(176,Y,32'b00000000000000000000000000000000,Z,1'b1,V,1'b0,N,1'b0);
  #10;

  //CASE: 177
  FN=6'b000111;
  A=32'b00010010001101000101011001111000;
  B=32'b00010010001101000101011001111000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(177,Y,32'b00000000000000000000000000000001,Z,1'b1,V,1'b0,N,1'b0);
  #10;

  //CASE: 178
  FN=6'b000011;
  A=32'b10000000000000000000000000000000;
  B=32'b00000000000000000000000000000001;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(178,Y,32'b00000000000000000000000000000000,Z,1'b0,V,1'b1,N,1'b0);
  #10;

  //CASE: 179
  FN=6'b000101;
  A=32'b10000000000000000000000000000000;
  B=32'b00000000000000000000000000000001;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(179,Y,32'b00000000000000000000000000000001,Z,1'b0,V,1'b1,N,1'b0);
  #10;

  //CASE: 180
  FN=6'b000111;
  A=32'b10000000000000000000000000000000;
  B=32'b00000000000000000000000000000001;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(180,Y,32'b00000000000000000000000000000001,Z,1'b0,V,1'b1,N,1'b0);
  #10;

  //CASE: 181
  FN=6'b000011;
  A=32'b11011110101011011011111011101111;
  B=32'b00000000000000000000000000000101;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(181,Y,32'b00000000000000000000000000000000,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 182
  FN=6'b000101;
  A=32'b11011110101011011011111011101111;
  B=32'b00000000000000000000000000000101;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(182,Y,32'b00000000000000000000000000000001,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 183
  FN=6'b000111;
  A=32'b11011110101011011011111011101111;
  B=32'b00000000000000000000000000000101;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(183,Y,32'b00000000000000000000000000000001,Z,1'b0,V,1'b0,N,1'b1);
  #10;

  //CASE: 184
  FN=6'b000011;
  A=32'b01111111111111111111111111111111;
  B=32'b11111111111111111111111111111111;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(184,Y,32'b00000000000000000000000000000000,Z,1'b0,V,1'b1,N,1'b1);
  #10;

  //CASE: 185
  FN=6'b000101;
  A=32'b01111111111111111111111111111111;
  B=32'b11111111111111111111111111111111;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(185,Y,32'b00000000000000000000000000000000,Z,1'b0,V,1'b1,N,1'b1);
  #10;

  //CASE: 186
  FN=6'b000111;
  A=32'b01111111111111111111111111111111;
  B=32'b11111111111111111111111111111111;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(186,Y,32'b00000000000000000000000000000000,Z,1'b0,V,1'b1,N,1'b1);
  #10;


  if(weAreOk) $display("TEST OK\n\nPassed");


  end

endmodule