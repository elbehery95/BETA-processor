`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Abdelrahman Elbehery
//
// Create Date:   00:32:16 02/10/2017
// Design Name:   BOOL
// Module Name:   F:/Self learning/FPGA/Projects/BETA_ISE/TB_BOOL.v
// Project Name:  BETA_ISE
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: BOOL
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module TB_BOOL;
  reg CLK=0;
  integer weAreOk=1;

  task PRINT;
    input integer CN;
    input [31:0] Y;
    input [31:0] ExY;
    if( Y!=ExY ) begin
    $display("Error in case: %d\nY: %b\nExpected: %b\n",CN,Y,ExY);
    weAreOk=0;
    end
  endtask

  reg [3:0] BFN;
  reg [31:0] A;
  reg [31:0] B;
  wire [31:0] Y;

  BOOL uut(.BFN(BFN),.A(A),.B(B),.Y(Y));



initial begin
  //CASE: 1
  BFN=4'b0000;
  A=32'b11111111000000001111111100000000;
  B=32'b11111111111111110000000000000000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(1,Y,32'b00000000000000000000000000000000);
  #10;

  //CASE: 2
  BFN=4'b0001;
  A=32'b11111111000000001111111100000000;
  B=32'b11111111111111110000000000000000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(2,Y,32'b00000000000000000000000011111111);
  #10;

  //CASE: 3
  BFN=4'b0010;
  A=32'b11111111000000001111111100000000;
  B=32'b11111111111111110000000000000000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(3,Y,32'b00000000000000001111111100000000);
  #10;

  //CASE: 4
  BFN=4'b0011;
  A=32'b11111111000000001111111100000000;
  B=32'b11111111111111110000000000000000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(4,Y,32'b00000000000000001111111111111111);
  #10;

  //CASE: 5
  BFN=4'b0100;
  A=32'b11111111000000001111111100000000;
  B=32'b11111111111111110000000000000000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(5,Y,32'b00000000111111110000000000000000);
  #10;

  //CASE: 6
  BFN=4'b0101;
  A=32'b11111111000000001111111100000000;
  B=32'b11111111111111110000000000000000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(6,Y,32'b00000000111111110000000011111111);
  #10;

  //CASE: 7
  BFN=4'b0110;
  A=32'b11111111000000001111111100000000;
  B=32'b11111111111111110000000000000000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(7,Y,32'b00000000111111111111111100000000);
  #10;

  //CASE: 8
  BFN=4'b0111;
  A=32'b11111111000000001111111100000000;
  B=32'b11111111111111110000000000000000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(8,Y,32'b00000000111111111111111111111111);
  #10;

  //CASE: 9
  BFN=4'b1000;
  A=32'b11111111000000001111111100000000;
  B=32'b11111111111111110000000000000000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(9,Y,32'b11111111000000000000000000000000);
  #10;

  //CASE: 10
  BFN=4'b1001;
  A=32'b11111111000000001111111100000000;
  B=32'b11111111111111110000000000000000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(10,Y,32'b11111111000000000000000011111111);
  #10;

  //CASE: 11
  BFN=4'b1010;
  A=32'b11111111000000001111111100000000;
  B=32'b11111111111111110000000000000000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(11,Y,32'b11111111000000001111111100000000);
  #10;

  //CASE: 12
  BFN=4'b1011;
  A=32'b11111111000000001111111100000000;
  B=32'b11111111111111110000000000000000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(12,Y,32'b11111111000000001111111111111111);
  #10;

  //CASE: 13
  BFN=4'b1100;
  A=32'b11111111000000001111111100000000;
  B=32'b11111111111111110000000000000000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(13,Y,32'b11111111111111110000000000000000);
  #10;

  //CASE: 14
  BFN=4'b1101;
  A=32'b11111111000000001111111100000000;
  B=32'b11111111111111110000000000000000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(14,Y,32'b11111111111111110000000011111111);
  #10;

  //CASE: 15
  BFN=4'b1110;
  A=32'b11111111000000001111111100000000;
  B=32'b11111111111111110000000000000000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(15,Y,32'b11111111111111111111111100000000);
  #10;

  //CASE: 16
  BFN=4'b1111;
  A=32'b11111111000000001111111100000000;
  B=32'b11111111111111110000000000000000;
  #1;
  CLK=1;
  #10;
  CLK=0;
  PRINT(16,Y,32'b11111111111111111111111111111111);
  #10;


  if(weAreOk) $display("TEST OK\n\nPassed");


  end

endmodule